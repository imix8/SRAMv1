* SPICE NETLIST
***************************************

.SUBCKT SRAMColumnNoCap !BL gnd! BL vdd! WL15 WL14 WL13 WL12 WL11 WL10 WL9 WL8 WL7 WL6 WL5 WL4 WL3 WL2 WL1 WL0
+ clk
** N=53 EP=21 IP=0 FDC=99
M0 3 WL15 !BL gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=1.79375e-14 AS=1.79375e-14 PD=5.55e-07 PS=5.55e-07 $X=2695 $Y=2665 $D=1
M1 4 WL14 !BL gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=1.79375e-14 AS=1.79375e-14 PD=5.55e-07 PS=5.55e-07 $X=2695 $Y=5125 $D=1
M2 5 WL13 !BL gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=1.79375e-14 AS=1.79375e-14 PD=5.55e-07 PS=5.55e-07 $X=2695 $Y=7610 $D=1
M3 6 WL12 !BL gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=1.79375e-14 AS=1.79375e-14 PD=5.55e-07 PS=5.55e-07 $X=2695 $Y=10070 $D=1
M4 7 WL11 !BL gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=1.79375e-14 AS=1.79375e-14 PD=5.55e-07 PS=5.55e-07 $X=2695 $Y=12530 $D=1
M5 8 WL10 !BL gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=1.79375e-14 AS=1.79375e-14 PD=5.55e-07 PS=5.55e-07 $X=2695 $Y=14990 $D=1
M6 9 WL9 !BL gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=1.79375e-14 AS=1.79375e-14 PD=5.55e-07 PS=5.55e-07 $X=2695 $Y=17475 $D=1
M7 10 WL8 !BL gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=1.79375e-14 AS=1.79375e-14 PD=5.55e-07 PS=5.55e-07 $X=2695 $Y=19935 $D=1
M8 11 WL7 !BL gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=1.79375e-14 AS=1.79375e-14 PD=5.55e-07 PS=5.55e-07 $X=2695 $Y=22395 $D=1
M9 12 WL6 !BL gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=1.79375e-14 AS=1.79375e-14 PD=5.55e-07 PS=5.55e-07 $X=2695 $Y=24855 $D=1
M10 13 WL5 !BL gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=1.79375e-14 AS=1.79375e-14 PD=5.55e-07 PS=5.55e-07 $X=2695 $Y=27340 $D=1
M11 14 WL4 !BL gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=1.79375e-14 AS=1.79375e-14 PD=5.55e-07 PS=5.55e-07 $X=2695 $Y=29800 $D=1
M12 15 WL3 !BL gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=1.79375e-14 AS=1.79375e-14 PD=5.55e-07 PS=5.55e-07 $X=2695 $Y=32260 $D=1
M13 16 WL2 !BL gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=1.79375e-14 AS=1.79375e-14 PD=5.55e-07 PS=5.55e-07 $X=2695 $Y=34720 $D=1
M14 17 WL1 !BL gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=1.79375e-14 AS=1.79375e-14 PD=5.55e-07 PS=5.55e-07 $X=2695 $Y=37205 $D=1
M15 18 WL0 !BL gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=1.79375e-14 AS=1.79375e-14 PD=5.55e-07 PS=5.55e-07 $X=2695 $Y=39665 $D=1
M16 20 3 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=2.05e-14 AS=2.05e-14 PD=6.05e-07 PS=6.05e-07 $X=3390 $Y=2645 $D=1
M17 21 4 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=2.05e-14 AS=2.05e-14 PD=6.05e-07 PS=6.05e-07 $X=3390 $Y=5105 $D=1
M18 22 5 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=2.05e-14 AS=2.05e-14 PD=6.05e-07 PS=6.05e-07 $X=3390 $Y=7590 $D=1
M19 23 6 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=2.05e-14 AS=2.05e-14 PD=6.05e-07 PS=6.05e-07 $X=3390 $Y=10050 $D=1
M20 24 7 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=2.05e-14 AS=2.05e-14 PD=6.05e-07 PS=6.05e-07 $X=3390 $Y=12510 $D=1
M21 25 8 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=2.05e-14 AS=2.05e-14 PD=6.05e-07 PS=6.05e-07 $X=3390 $Y=14970 $D=1
M22 26 9 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=2.05e-14 AS=2.05e-14 PD=6.05e-07 PS=6.05e-07 $X=3390 $Y=17455 $D=1
M23 27 10 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=2.05e-14 AS=2.05e-14 PD=6.05e-07 PS=6.05e-07 $X=3390 $Y=19915 $D=1
M24 28 11 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=2.05e-14 AS=2.05e-14 PD=6.05e-07 PS=6.05e-07 $X=3390 $Y=22375 $D=1
M25 29 12 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=2.05e-14 AS=2.05e-14 PD=6.05e-07 PS=6.05e-07 $X=3390 $Y=24835 $D=1
M26 30 13 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=2.05e-14 AS=2.05e-14 PD=6.05e-07 PS=6.05e-07 $X=3390 $Y=27320 $D=1
M27 31 14 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=2.05e-14 AS=2.05e-14 PD=6.05e-07 PS=6.05e-07 $X=3390 $Y=29780 $D=1
M28 32 15 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=2.05e-14 AS=2.05e-14 PD=6.05e-07 PS=6.05e-07 $X=3390 $Y=32240 $D=1
M29 33 16 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=2.05e-14 AS=2.05e-14 PD=6.05e-07 PS=6.05e-07 $X=3390 $Y=34700 $D=1
M30 34 17 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=2.05e-14 AS=2.05e-14 PD=6.05e-07 PS=6.05e-07 $X=3390 $Y=37185 $D=1
M31 35 18 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=2.05e-14 AS=2.05e-14 PD=6.05e-07 PS=6.05e-07 $X=3390 $Y=39645 $D=1
M32 gnd! 20 3 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=2.05e-14 AS=2.05e-14 PD=6.05e-07 PS=6.05e-07 $X=4160 $Y=2645 $D=1
M33 gnd! 21 4 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=2.05e-14 AS=2.05e-14 PD=6.05e-07 PS=6.05e-07 $X=4160 $Y=5105 $D=1
M34 gnd! 22 5 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=2.05e-14 AS=2.05e-14 PD=6.05e-07 PS=6.05e-07 $X=4160 $Y=7590 $D=1
M35 gnd! 23 6 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=2.05e-14 AS=2.05e-14 PD=6.05e-07 PS=6.05e-07 $X=4160 $Y=10050 $D=1
M36 gnd! 24 7 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=2.05e-14 AS=2.05e-14 PD=6.05e-07 PS=6.05e-07 $X=4160 $Y=12510 $D=1
M37 gnd! 25 8 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=2.05e-14 AS=2.05e-14 PD=6.05e-07 PS=6.05e-07 $X=4160 $Y=14970 $D=1
M38 gnd! 26 9 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=2.05e-14 AS=2.05e-14 PD=6.05e-07 PS=6.05e-07 $X=4160 $Y=17455 $D=1
M39 gnd! 27 10 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=2.05e-14 AS=2.05e-14 PD=6.05e-07 PS=6.05e-07 $X=4160 $Y=19915 $D=1
M40 gnd! 28 11 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=2.05e-14 AS=2.05e-14 PD=6.05e-07 PS=6.05e-07 $X=4160 $Y=22375 $D=1
M41 gnd! 29 12 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=2.05e-14 AS=2.05e-14 PD=6.05e-07 PS=6.05e-07 $X=4160 $Y=24835 $D=1
M42 gnd! 30 13 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=2.05e-14 AS=2.05e-14 PD=6.05e-07 PS=6.05e-07 $X=4160 $Y=27320 $D=1
M43 gnd! 31 14 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=2.05e-14 AS=2.05e-14 PD=6.05e-07 PS=6.05e-07 $X=4160 $Y=29780 $D=1
M44 gnd! 32 15 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=2.05e-14 AS=2.05e-14 PD=6.05e-07 PS=6.05e-07 $X=4160 $Y=32240 $D=1
M45 gnd! 33 16 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=2.05e-14 AS=2.05e-14 PD=6.05e-07 PS=6.05e-07 $X=4160 $Y=34700 $D=1
M46 gnd! 34 17 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=2.05e-14 AS=2.05e-14 PD=6.05e-07 PS=6.05e-07 $X=4160 $Y=37185 $D=1
M47 gnd! 35 18 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=2.05e-14 AS=2.05e-14 PD=6.05e-07 PS=6.05e-07 $X=4160 $Y=39645 $D=1
M48 BL WL15 20 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=1.79375e-14 AS=1.79375e-14 PD=5.55e-07 PS=5.55e-07 $X=4840 $Y=2675 $D=1
M49 BL WL14 21 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=1.79375e-14 AS=1.79375e-14 PD=5.55e-07 PS=5.55e-07 $X=4840 $Y=5135 $D=1
M50 BL WL13 22 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=1.79375e-14 AS=1.79375e-14 PD=5.55e-07 PS=5.55e-07 $X=4840 $Y=7620 $D=1
M51 BL WL12 23 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=1.79375e-14 AS=1.79375e-14 PD=5.55e-07 PS=5.55e-07 $X=4840 $Y=10080 $D=1
M52 BL WL11 24 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=1.79375e-14 AS=1.79375e-14 PD=5.55e-07 PS=5.55e-07 $X=4840 $Y=12540 $D=1
M53 BL WL10 25 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=1.79375e-14 AS=1.79375e-14 PD=5.55e-07 PS=5.55e-07 $X=4840 $Y=15000 $D=1
M54 BL WL9 26 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=1.79375e-14 AS=1.79375e-14 PD=5.55e-07 PS=5.55e-07 $X=4840 $Y=17485 $D=1
M55 BL WL8 27 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=1.79375e-14 AS=1.79375e-14 PD=5.55e-07 PS=5.55e-07 $X=4840 $Y=19945 $D=1
M56 BL WL7 28 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=1.79375e-14 AS=1.79375e-14 PD=5.55e-07 PS=5.55e-07 $X=4840 $Y=22405 $D=1
M57 BL WL6 29 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=1.79375e-14 AS=1.79375e-14 PD=5.55e-07 PS=5.55e-07 $X=4840 $Y=24865 $D=1
M58 BL WL5 30 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=1.79375e-14 AS=1.79375e-14 PD=5.55e-07 PS=5.55e-07 $X=4840 $Y=27350 $D=1
M59 BL WL4 31 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=1.79375e-14 AS=1.79375e-14 PD=5.55e-07 PS=5.55e-07 $X=4840 $Y=29810 $D=1
M60 BL WL3 32 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=1.79375e-14 AS=1.79375e-14 PD=5.55e-07 PS=5.55e-07 $X=4840 $Y=32270 $D=1
M61 BL WL2 33 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=1.79375e-14 AS=1.79375e-14 PD=5.55e-07 PS=5.55e-07 $X=4840 $Y=34730 $D=1
M62 BL WL1 34 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=1.79375e-14 AS=1.79375e-14 PD=5.55e-07 PS=5.55e-07 $X=4840 $Y=37215 $D=1
M63 BL WL0 35 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=1.79375e-14 AS=1.79375e-14 PD=5.55e-07 PS=5.55e-07 $X=4840 $Y=39675 $D=1
M64 BL clk vdd! vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=2825 $Y=42100 $D=0
M65 20 3 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.025e-14 AS=1.025e-14 PD=4.05e-07 PS=4.05e-07 $X=3390 $Y=3825 $D=0
M66 21 4 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.025e-14 AS=1.025e-14 PD=4.05e-07 PS=4.05e-07 $X=3390 $Y=6285 $D=0
M67 22 5 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.025e-14 AS=1.025e-14 PD=4.05e-07 PS=4.05e-07 $X=3390 $Y=8770 $D=0
M68 23 6 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.025e-14 AS=1.025e-14 PD=4.05e-07 PS=4.05e-07 $X=3390 $Y=11230 $D=0
M69 24 7 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.025e-14 AS=1.025e-14 PD=4.05e-07 PS=4.05e-07 $X=3390 $Y=13690 $D=0
M70 25 8 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.025e-14 AS=1.025e-14 PD=4.05e-07 PS=4.05e-07 $X=3390 $Y=16150 $D=0
M71 26 9 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.025e-14 AS=1.025e-14 PD=4.05e-07 PS=4.05e-07 $X=3390 $Y=18635 $D=0
M72 27 10 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.025e-14 AS=1.025e-14 PD=4.05e-07 PS=4.05e-07 $X=3390 $Y=21095 $D=0
M73 28 11 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.025e-14 AS=1.025e-14 PD=4.05e-07 PS=4.05e-07 $X=3390 $Y=23555 $D=0
M74 29 12 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.025e-14 AS=1.025e-14 PD=4.05e-07 PS=4.05e-07 $X=3390 $Y=26015 $D=0
M75 30 13 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.025e-14 AS=1.025e-14 PD=4.05e-07 PS=4.05e-07 $X=3390 $Y=28500 $D=0
M76 31 14 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.025e-14 AS=1.025e-14 PD=4.05e-07 PS=4.05e-07 $X=3390 $Y=30960 $D=0
M77 32 15 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.025e-14 AS=1.025e-14 PD=4.05e-07 PS=4.05e-07 $X=3390 $Y=33420 $D=0
M78 33 16 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.025e-14 AS=1.025e-14 PD=4.05e-07 PS=4.05e-07 $X=3390 $Y=35880 $D=0
M79 34 17 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.025e-14 AS=1.025e-14 PD=4.05e-07 PS=4.05e-07 $X=3390 $Y=38365 $D=0
M80 35 18 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.025e-14 AS=1.025e-14 PD=4.05e-07 PS=4.05e-07 $X=3390 $Y=40825 $D=0
M81 !BL clk BL vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=3680 $Y=42100 $D=0
M82 vdd! 20 3 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.025e-14 AS=1.025e-14 PD=4.05e-07 PS=4.05e-07 $X=4160 $Y=3825 $D=0
M83 vdd! 21 4 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.025e-14 AS=1.025e-14 PD=4.05e-07 PS=4.05e-07 $X=4160 $Y=6285 $D=0
M84 vdd! 22 5 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.025e-14 AS=1.025e-14 PD=4.05e-07 PS=4.05e-07 $X=4160 $Y=8770 $D=0
M85 vdd! 23 6 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.025e-14 AS=1.025e-14 PD=4.05e-07 PS=4.05e-07 $X=4160 $Y=11230 $D=0
M86 vdd! 24 7 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.025e-14 AS=1.025e-14 PD=4.05e-07 PS=4.05e-07 $X=4160 $Y=13690 $D=0
M87 vdd! 25 8 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.025e-14 AS=1.025e-14 PD=4.05e-07 PS=4.05e-07 $X=4160 $Y=16150 $D=0
M88 vdd! 26 9 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.025e-14 AS=1.025e-14 PD=4.05e-07 PS=4.05e-07 $X=4160 $Y=18635 $D=0
M89 vdd! 27 10 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.025e-14 AS=1.025e-14 PD=4.05e-07 PS=4.05e-07 $X=4160 $Y=21095 $D=0
M90 vdd! 28 11 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.025e-14 AS=1.025e-14 PD=4.05e-07 PS=4.05e-07 $X=4160 $Y=23555 $D=0
M91 vdd! 29 12 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.025e-14 AS=1.025e-14 PD=4.05e-07 PS=4.05e-07 $X=4160 $Y=26015 $D=0
M92 vdd! 30 13 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.025e-14 AS=1.025e-14 PD=4.05e-07 PS=4.05e-07 $X=4160 $Y=28500 $D=0
M93 vdd! 31 14 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.025e-14 AS=1.025e-14 PD=4.05e-07 PS=4.05e-07 $X=4160 $Y=30960 $D=0
M94 vdd! 32 15 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.025e-14 AS=1.025e-14 PD=4.05e-07 PS=4.05e-07 $X=4160 $Y=33420 $D=0
M95 vdd! 33 16 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.025e-14 AS=1.025e-14 PD=4.05e-07 PS=4.05e-07 $X=4160 $Y=35880 $D=0
M96 vdd! 34 17 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.025e-14 AS=1.025e-14 PD=4.05e-07 PS=4.05e-07 $X=4160 $Y=38365 $D=0
M97 vdd! 35 18 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.025e-14 AS=1.025e-14 PD=4.05e-07 PS=4.05e-07 $X=4160 $Y=40825 $D=0
M98 vdd! clk !BL vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=4545 $Y=42100 $D=0
.ENDS
***************************************
