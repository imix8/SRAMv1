* SPICE NETLIST
***************************************

.SUBCKT SRAMArray gnd! !BL0 BL0 !BL1 BL1 !BL2 BL2 !BL3 BL3 !BL4 BL4 !BL5 BL5 !BL6 BL6 !BL7 BL7 !BL8 BL8 !BL9
+ BL9 !BL10 BL10 !BL11 BL11 !BL12 BL12 !BL13 BL13 !BL14 BL14 !BL15 BL15 !BL16 BL16 !BL17 BL17 !BL18 BL18 !BL19
+ BL19 !BL20 BL20 !BL21 BL21 !BL22 BL22 !BL23 BL23 !BL24 BL24 !BL25 BL25 !BL26 BL26 !BL27 BL27 !BL28 BL28 !BL29
+ BL29 !BL30 BL30 !BL31 BL31 WL15 WL14 WL13 WL12 WL11 WL10 WL9 WL8 WL7 WL6 WL5 WL4 WL3 WL2 WL1
+ WL0 clk vdd!
** N=1107 EP=83 IP=0 FDC=3168
M0 82 WL15 !BL0 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=1175 $Y=1085 $D=1
M1 83 WL14 !BL0 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=1175 $Y=4575 $D=1
M2 84 WL13 !BL0 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=1175 $Y=8065 $D=1
M3 85 WL12 !BL0 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=1175 $Y=11555 $D=1
M4 86 WL11 !BL0 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=1175 $Y=15045 $D=1
M5 87 WL10 !BL0 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=1175 $Y=18535 $D=1
M6 88 WL9 !BL0 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=1175 $Y=22025 $D=1
M7 89 WL8 !BL0 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=1175 $Y=25515 $D=1
M8 90 WL7 !BL0 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=1175 $Y=29005 $D=1
M9 91 WL6 !BL0 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=1175 $Y=32495 $D=1
M10 92 WL5 !BL0 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=1175 $Y=35985 $D=1
M11 93 WL4 !BL0 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=1175 $Y=39475 $D=1
M12 94 WL3 !BL0 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=1175 $Y=42965 $D=1
M13 95 WL2 !BL0 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=1175 $Y=46455 $D=1
M14 96 WL1 !BL0 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=1175 $Y=49945 $D=1
M15 97 WL0 !BL0 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=1175 $Y=53435 $D=1
M16 gnd! 99 82 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=1900 $Y=1330 $D=1
M17 gnd! 100 83 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=1900 $Y=4820 $D=1
M18 gnd! 101 84 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=1900 $Y=8310 $D=1
M19 gnd! 102 85 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=1900 $Y=11800 $D=1
M20 gnd! 103 86 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=1900 $Y=15290 $D=1
M21 gnd! 104 87 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=1900 $Y=18780 $D=1
M22 gnd! 105 88 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=1900 $Y=22270 $D=1
M23 gnd! 106 89 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=1900 $Y=25760 $D=1
M24 gnd! 107 90 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=1900 $Y=29250 $D=1
M25 gnd! 108 91 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=1900 $Y=32740 $D=1
M26 gnd! 109 92 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=1900 $Y=36230 $D=1
M27 gnd! 110 93 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=1900 $Y=39720 $D=1
M28 gnd! 111 94 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=1900 $Y=43210 $D=1
M29 gnd! 112 95 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=1900 $Y=46700 $D=1
M30 gnd! 113 96 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=1900 $Y=50190 $D=1
M31 gnd! 114 97 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=1900 $Y=53680 $D=1
M32 99 82 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=2490 $Y=1330 $D=1
M33 100 83 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=2490 $Y=4820 $D=1
M34 101 84 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=2490 $Y=8310 $D=1
M35 102 85 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=2490 $Y=11800 $D=1
M36 103 86 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=2490 $Y=15290 $D=1
M37 104 87 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=2490 $Y=18780 $D=1
M38 105 88 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=2490 $Y=22270 $D=1
M39 106 89 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=2490 $Y=25760 $D=1
M40 107 90 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=2490 $Y=29250 $D=1
M41 108 91 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=2490 $Y=32740 $D=1
M42 109 92 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=2490 $Y=36230 $D=1
M43 110 93 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=2490 $Y=39720 $D=1
M44 111 94 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=2490 $Y=43210 $D=1
M45 112 95 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=2490 $Y=46700 $D=1
M46 113 96 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=2490 $Y=50190 $D=1
M47 114 97 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=2490 $Y=53680 $D=1
M48 99 WL15 BL0 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=2930 $Y=1085 $D=1
M49 100 WL14 BL0 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=2930 $Y=4575 $D=1
M50 101 WL13 BL0 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=2930 $Y=8065 $D=1
M51 102 WL12 BL0 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=2930 $Y=11555 $D=1
M52 103 WL11 BL0 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=2930 $Y=15045 $D=1
M53 104 WL10 BL0 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=2930 $Y=18535 $D=1
M54 105 WL9 BL0 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=2930 $Y=22025 $D=1
M55 106 WL8 BL0 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=2930 $Y=25515 $D=1
M56 107 WL7 BL0 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=2930 $Y=29005 $D=1
M57 108 WL6 BL0 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=2930 $Y=32495 $D=1
M58 109 WL5 BL0 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=2930 $Y=35985 $D=1
M59 110 WL4 BL0 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=2930 $Y=39475 $D=1
M60 111 WL3 BL0 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=2930 $Y=42965 $D=1
M61 112 WL2 BL0 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=2930 $Y=46455 $D=1
M62 113 WL1 BL0 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=2930 $Y=49945 $D=1
M63 114 WL0 BL0 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=2930 $Y=53435 $D=1
M64 115 WL15 !BL1 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=4280 $Y=1085 $D=1
M65 116 WL14 !BL1 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=4280 $Y=4575 $D=1
M66 117 WL13 !BL1 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=4280 $Y=8065 $D=1
M67 118 WL12 !BL1 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=4280 $Y=11555 $D=1
M68 119 WL11 !BL1 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=4280 $Y=15045 $D=1
M69 120 WL10 !BL1 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=4280 $Y=18535 $D=1
M70 121 WL9 !BL1 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=4280 $Y=22025 $D=1
M71 122 WL8 !BL1 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=4280 $Y=25515 $D=1
M72 123 WL7 !BL1 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=4280 $Y=29005 $D=1
M73 124 WL6 !BL1 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=4280 $Y=32495 $D=1
M74 125 WL5 !BL1 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=4280 $Y=35985 $D=1
M75 126 WL4 !BL1 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=4280 $Y=39475 $D=1
M76 127 WL3 !BL1 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=4280 $Y=42965 $D=1
M77 128 WL2 !BL1 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=4280 $Y=46455 $D=1
M78 129 WL1 !BL1 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=4280 $Y=49945 $D=1
M79 130 WL0 !BL1 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=4280 $Y=53435 $D=1
M80 gnd! 131 115 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=5005 $Y=1330 $D=1
M81 gnd! 132 116 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=5005 $Y=4820 $D=1
M82 gnd! 133 117 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=5005 $Y=8310 $D=1
M83 gnd! 134 118 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=5005 $Y=11800 $D=1
M84 gnd! 135 119 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=5005 $Y=15290 $D=1
M85 gnd! 136 120 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=5005 $Y=18780 $D=1
M86 gnd! 137 121 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=5005 $Y=22270 $D=1
M87 gnd! 138 122 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=5005 $Y=25760 $D=1
M88 gnd! 139 123 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=5005 $Y=29250 $D=1
M89 gnd! 140 124 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=5005 $Y=32740 $D=1
M90 gnd! 141 125 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=5005 $Y=36230 $D=1
M91 gnd! 142 126 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=5005 $Y=39720 $D=1
M92 gnd! 143 127 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=5005 $Y=43210 $D=1
M93 gnd! 144 128 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=5005 $Y=46700 $D=1
M94 gnd! 145 129 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=5005 $Y=50190 $D=1
M95 gnd! 146 130 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=5005 $Y=53680 $D=1
M96 131 115 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=5595 $Y=1330 $D=1
M97 132 116 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=5595 $Y=4820 $D=1
M98 133 117 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=5595 $Y=8310 $D=1
M99 134 118 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=5595 $Y=11800 $D=1
M100 135 119 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=5595 $Y=15290 $D=1
M101 136 120 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=5595 $Y=18780 $D=1
M102 137 121 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=5595 $Y=22270 $D=1
M103 138 122 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=5595 $Y=25760 $D=1
M104 139 123 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=5595 $Y=29250 $D=1
M105 140 124 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=5595 $Y=32740 $D=1
M106 141 125 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=5595 $Y=36230 $D=1
M107 142 126 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=5595 $Y=39720 $D=1
M108 143 127 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=5595 $Y=43210 $D=1
M109 144 128 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=5595 $Y=46700 $D=1
M110 145 129 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=5595 $Y=50190 $D=1
M111 146 130 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=5595 $Y=53680 $D=1
M112 131 WL15 BL1 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=6035 $Y=1085 $D=1
M113 132 WL14 BL1 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=6035 $Y=4575 $D=1
M114 133 WL13 BL1 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=6035 $Y=8065 $D=1
M115 134 WL12 BL1 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=6035 $Y=11555 $D=1
M116 135 WL11 BL1 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=6035 $Y=15045 $D=1
M117 136 WL10 BL1 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=6035 $Y=18535 $D=1
M118 137 WL9 BL1 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=6035 $Y=22025 $D=1
M119 138 WL8 BL1 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=6035 $Y=25515 $D=1
M120 139 WL7 BL1 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=6035 $Y=29005 $D=1
M121 140 WL6 BL1 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=6035 $Y=32495 $D=1
M122 141 WL5 BL1 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=6035 $Y=35985 $D=1
M123 142 WL4 BL1 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=6035 $Y=39475 $D=1
M124 143 WL3 BL1 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=6035 $Y=42965 $D=1
M125 144 WL2 BL1 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=6035 $Y=46455 $D=1
M126 145 WL1 BL1 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=6035 $Y=49945 $D=1
M127 146 WL0 BL1 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=6035 $Y=53435 $D=1
M128 147 WL15 !BL2 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=7385 $Y=1085 $D=1
M129 148 WL14 !BL2 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=7385 $Y=4575 $D=1
M130 149 WL13 !BL2 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=7385 $Y=8065 $D=1
M131 150 WL12 !BL2 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=7385 $Y=11555 $D=1
M132 151 WL11 !BL2 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=7385 $Y=15045 $D=1
M133 152 WL10 !BL2 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=7385 $Y=18535 $D=1
M134 153 WL9 !BL2 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=7385 $Y=22025 $D=1
M135 154 WL8 !BL2 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=7385 $Y=25515 $D=1
M136 155 WL7 !BL2 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=7385 $Y=29005 $D=1
M137 156 WL6 !BL2 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=7385 $Y=32495 $D=1
M138 157 WL5 !BL2 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=7385 $Y=35985 $D=1
M139 158 WL4 !BL2 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=7385 $Y=39475 $D=1
M140 159 WL3 !BL2 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=7385 $Y=42965 $D=1
M141 160 WL2 !BL2 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=7385 $Y=46455 $D=1
M142 161 WL1 !BL2 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=7385 $Y=49945 $D=1
M143 162 WL0 !BL2 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=7385 $Y=53435 $D=1
M144 gnd! 163 147 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=8110 $Y=1330 $D=1
M145 gnd! 164 148 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=8110 $Y=4820 $D=1
M146 gnd! 165 149 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=8110 $Y=8310 $D=1
M147 gnd! 166 150 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=8110 $Y=11800 $D=1
M148 gnd! 167 151 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=8110 $Y=15290 $D=1
M149 gnd! 168 152 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=8110 $Y=18780 $D=1
M150 gnd! 169 153 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=8110 $Y=22270 $D=1
M151 gnd! 170 154 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=8110 $Y=25760 $D=1
M152 gnd! 171 155 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=8110 $Y=29250 $D=1
M153 gnd! 172 156 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=8110 $Y=32740 $D=1
M154 gnd! 173 157 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=8110 $Y=36230 $D=1
M155 gnd! 174 158 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=8110 $Y=39720 $D=1
M156 gnd! 175 159 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=8110 $Y=43210 $D=1
M157 gnd! 176 160 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=8110 $Y=46700 $D=1
M158 gnd! 177 161 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=8110 $Y=50190 $D=1
M159 gnd! 178 162 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=8110 $Y=53680 $D=1
M160 163 147 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=8700 $Y=1330 $D=1
M161 164 148 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=8700 $Y=4820 $D=1
M162 165 149 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=8700 $Y=8310 $D=1
M163 166 150 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=8700 $Y=11800 $D=1
M164 167 151 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=8700 $Y=15290 $D=1
M165 168 152 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=8700 $Y=18780 $D=1
M166 169 153 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=8700 $Y=22270 $D=1
M167 170 154 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=8700 $Y=25760 $D=1
M168 171 155 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=8700 $Y=29250 $D=1
M169 172 156 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=8700 $Y=32740 $D=1
M170 173 157 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=8700 $Y=36230 $D=1
M171 174 158 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=8700 $Y=39720 $D=1
M172 175 159 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=8700 $Y=43210 $D=1
M173 176 160 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=8700 $Y=46700 $D=1
M174 177 161 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=8700 $Y=50190 $D=1
M175 178 162 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=8700 $Y=53680 $D=1
M176 163 WL15 BL2 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=9140 $Y=1085 $D=1
M177 164 WL14 BL2 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=9140 $Y=4575 $D=1
M178 165 WL13 BL2 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=9140 $Y=8065 $D=1
M179 166 WL12 BL2 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=9140 $Y=11555 $D=1
M180 167 WL11 BL2 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=9140 $Y=15045 $D=1
M181 168 WL10 BL2 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=9140 $Y=18535 $D=1
M182 169 WL9 BL2 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=9140 $Y=22025 $D=1
M183 170 WL8 BL2 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=9140 $Y=25515 $D=1
M184 171 WL7 BL2 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=9140 $Y=29005 $D=1
M185 172 WL6 BL2 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=9140 $Y=32495 $D=1
M186 173 WL5 BL2 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=9140 $Y=35985 $D=1
M187 174 WL4 BL2 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=9140 $Y=39475 $D=1
M188 175 WL3 BL2 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=9140 $Y=42965 $D=1
M189 176 WL2 BL2 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=9140 $Y=46455 $D=1
M190 177 WL1 BL2 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=9140 $Y=49945 $D=1
M191 178 WL0 BL2 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=9140 $Y=53435 $D=1
M192 179 WL15 !BL3 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=10490 $Y=1085 $D=1
M193 180 WL14 !BL3 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=10490 $Y=4575 $D=1
M194 181 WL13 !BL3 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=10490 $Y=8065 $D=1
M195 182 WL12 !BL3 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=10490 $Y=11555 $D=1
M196 183 WL11 !BL3 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=10490 $Y=15045 $D=1
M197 184 WL10 !BL3 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=10490 $Y=18535 $D=1
M198 185 WL9 !BL3 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=10490 $Y=22025 $D=1
M199 186 WL8 !BL3 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=10490 $Y=25515 $D=1
M200 187 WL7 !BL3 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=10490 $Y=29005 $D=1
M201 188 WL6 !BL3 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=10490 $Y=32495 $D=1
M202 189 WL5 !BL3 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=10490 $Y=35985 $D=1
M203 190 WL4 !BL3 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=10490 $Y=39475 $D=1
M204 191 WL3 !BL3 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=10490 $Y=42965 $D=1
M205 192 WL2 !BL3 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=10490 $Y=46455 $D=1
M206 193 WL1 !BL3 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=10490 $Y=49945 $D=1
M207 194 WL0 !BL3 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=10490 $Y=53435 $D=1
M208 gnd! 195 179 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=11215 $Y=1330 $D=1
M209 gnd! 196 180 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=11215 $Y=4820 $D=1
M210 gnd! 197 181 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=11215 $Y=8310 $D=1
M211 gnd! 198 182 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=11215 $Y=11800 $D=1
M212 gnd! 199 183 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=11215 $Y=15290 $D=1
M213 gnd! 200 184 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=11215 $Y=18780 $D=1
M214 gnd! 201 185 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=11215 $Y=22270 $D=1
M215 gnd! 202 186 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=11215 $Y=25760 $D=1
M216 gnd! 203 187 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=11215 $Y=29250 $D=1
M217 gnd! 204 188 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=11215 $Y=32740 $D=1
M218 gnd! 205 189 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=11215 $Y=36230 $D=1
M219 gnd! 206 190 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=11215 $Y=39720 $D=1
M220 gnd! 207 191 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=11215 $Y=43210 $D=1
M221 gnd! 208 192 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=11215 $Y=46700 $D=1
M222 gnd! 209 193 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=11215 $Y=50190 $D=1
M223 gnd! 210 194 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=11215 $Y=53680 $D=1
M224 195 179 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=11805 $Y=1330 $D=1
M225 196 180 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=11805 $Y=4820 $D=1
M226 197 181 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=11805 $Y=8310 $D=1
M227 198 182 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=11805 $Y=11800 $D=1
M228 199 183 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=11805 $Y=15290 $D=1
M229 200 184 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=11805 $Y=18780 $D=1
M230 201 185 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=11805 $Y=22270 $D=1
M231 202 186 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=11805 $Y=25760 $D=1
M232 203 187 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=11805 $Y=29250 $D=1
M233 204 188 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=11805 $Y=32740 $D=1
M234 205 189 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=11805 $Y=36230 $D=1
M235 206 190 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=11805 $Y=39720 $D=1
M236 207 191 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=11805 $Y=43210 $D=1
M237 208 192 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=11805 $Y=46700 $D=1
M238 209 193 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=11805 $Y=50190 $D=1
M239 210 194 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=11805 $Y=53680 $D=1
M240 195 WL15 BL3 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=12245 $Y=1085 $D=1
M241 196 WL14 BL3 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=12245 $Y=4575 $D=1
M242 197 WL13 BL3 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=12245 $Y=8065 $D=1
M243 198 WL12 BL3 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=12245 $Y=11555 $D=1
M244 199 WL11 BL3 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=12245 $Y=15045 $D=1
M245 200 WL10 BL3 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=12245 $Y=18535 $D=1
M246 201 WL9 BL3 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=12245 $Y=22025 $D=1
M247 202 WL8 BL3 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=12245 $Y=25515 $D=1
M248 203 WL7 BL3 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=12245 $Y=29005 $D=1
M249 204 WL6 BL3 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=12245 $Y=32495 $D=1
M250 205 WL5 BL3 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=12245 $Y=35985 $D=1
M251 206 WL4 BL3 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=12245 $Y=39475 $D=1
M252 207 WL3 BL3 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=12245 $Y=42965 $D=1
M253 208 WL2 BL3 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=12245 $Y=46455 $D=1
M254 209 WL1 BL3 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=12245 $Y=49945 $D=1
M255 210 WL0 BL3 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=12245 $Y=53435 $D=1
M256 211 WL15 !BL4 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=13595 $Y=1085 $D=1
M257 212 WL14 !BL4 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=13595 $Y=4575 $D=1
M258 213 WL13 !BL4 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=13595 $Y=8065 $D=1
M259 214 WL12 !BL4 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=13595 $Y=11555 $D=1
M260 215 WL11 !BL4 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=13595 $Y=15045 $D=1
M261 216 WL10 !BL4 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=13595 $Y=18535 $D=1
M262 217 WL9 !BL4 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=13595 $Y=22025 $D=1
M263 218 WL8 !BL4 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=13595 $Y=25515 $D=1
M264 219 WL7 !BL4 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=13595 $Y=29005 $D=1
M265 220 WL6 !BL4 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=13595 $Y=32495 $D=1
M266 221 WL5 !BL4 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=13595 $Y=35985 $D=1
M267 222 WL4 !BL4 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=13595 $Y=39475 $D=1
M268 223 WL3 !BL4 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=13595 $Y=42965 $D=1
M269 224 WL2 !BL4 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=13595 $Y=46455 $D=1
M270 225 WL1 !BL4 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=13595 $Y=49945 $D=1
M271 226 WL0 !BL4 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=13595 $Y=53435 $D=1
M272 gnd! 227 211 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=14320 $Y=1330 $D=1
M273 gnd! 228 212 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=14320 $Y=4820 $D=1
M274 gnd! 229 213 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=14320 $Y=8310 $D=1
M275 gnd! 230 214 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=14320 $Y=11800 $D=1
M276 gnd! 231 215 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=14320 $Y=15290 $D=1
M277 gnd! 232 216 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=14320 $Y=18780 $D=1
M278 gnd! 233 217 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=14320 $Y=22270 $D=1
M279 gnd! 234 218 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=14320 $Y=25760 $D=1
M280 gnd! 235 219 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=14320 $Y=29250 $D=1
M281 gnd! 236 220 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=14320 $Y=32740 $D=1
M282 gnd! 237 221 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=14320 $Y=36230 $D=1
M283 gnd! 238 222 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=14320 $Y=39720 $D=1
M284 gnd! 239 223 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=14320 $Y=43210 $D=1
M285 gnd! 240 224 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=14320 $Y=46700 $D=1
M286 gnd! 241 225 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=14320 $Y=50190 $D=1
M287 gnd! 242 226 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=14320 $Y=53680 $D=1
M288 227 211 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=14910 $Y=1330 $D=1
M289 228 212 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=14910 $Y=4820 $D=1
M290 229 213 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=14910 $Y=8310 $D=1
M291 230 214 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=14910 $Y=11800 $D=1
M292 231 215 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=14910 $Y=15290 $D=1
M293 232 216 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=14910 $Y=18780 $D=1
M294 233 217 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=14910 $Y=22270 $D=1
M295 234 218 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=14910 $Y=25760 $D=1
M296 235 219 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=14910 $Y=29250 $D=1
M297 236 220 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=14910 $Y=32740 $D=1
M298 237 221 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=14910 $Y=36230 $D=1
M299 238 222 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=14910 $Y=39720 $D=1
M300 239 223 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=14910 $Y=43210 $D=1
M301 240 224 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=14910 $Y=46700 $D=1
M302 241 225 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=14910 $Y=50190 $D=1
M303 242 226 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=14910 $Y=53680 $D=1
M304 227 WL15 BL4 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=15350 $Y=1085 $D=1
M305 228 WL14 BL4 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=15350 $Y=4575 $D=1
M306 229 WL13 BL4 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=15350 $Y=8065 $D=1
M307 230 WL12 BL4 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=15350 $Y=11555 $D=1
M308 231 WL11 BL4 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=15350 $Y=15045 $D=1
M309 232 WL10 BL4 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=15350 $Y=18535 $D=1
M310 233 WL9 BL4 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=15350 $Y=22025 $D=1
M311 234 WL8 BL4 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=15350 $Y=25515 $D=1
M312 235 WL7 BL4 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=15350 $Y=29005 $D=1
M313 236 WL6 BL4 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=15350 $Y=32495 $D=1
M314 237 WL5 BL4 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=15350 $Y=35985 $D=1
M315 238 WL4 BL4 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=15350 $Y=39475 $D=1
M316 239 WL3 BL4 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=15350 $Y=42965 $D=1
M317 240 WL2 BL4 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=15350 $Y=46455 $D=1
M318 241 WL1 BL4 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=15350 $Y=49945 $D=1
M319 242 WL0 BL4 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=15350 $Y=53435 $D=1
M320 243 WL15 !BL5 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=16700 $Y=1085 $D=1
M321 244 WL14 !BL5 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=16700 $Y=4575 $D=1
M322 245 WL13 !BL5 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=16700 $Y=8065 $D=1
M323 246 WL12 !BL5 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=16700 $Y=11555 $D=1
M324 247 WL11 !BL5 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=16700 $Y=15045 $D=1
M325 248 WL10 !BL5 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=16700 $Y=18535 $D=1
M326 249 WL9 !BL5 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=16700 $Y=22025 $D=1
M327 250 WL8 !BL5 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=16700 $Y=25515 $D=1
M328 251 WL7 !BL5 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=16700 $Y=29005 $D=1
M329 252 WL6 !BL5 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=16700 $Y=32495 $D=1
M330 253 WL5 !BL5 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=16700 $Y=35985 $D=1
M331 254 WL4 !BL5 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=16700 $Y=39475 $D=1
M332 255 WL3 !BL5 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=16700 $Y=42965 $D=1
M333 256 WL2 !BL5 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=16700 $Y=46455 $D=1
M334 257 WL1 !BL5 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=16700 $Y=49945 $D=1
M335 258 WL0 !BL5 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=16700 $Y=53435 $D=1
M336 gnd! 259 243 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=17425 $Y=1330 $D=1
M337 gnd! 260 244 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=17425 $Y=4820 $D=1
M338 gnd! 261 245 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=17425 $Y=8310 $D=1
M339 gnd! 262 246 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=17425 $Y=11800 $D=1
M340 gnd! 263 247 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=17425 $Y=15290 $D=1
M341 gnd! 264 248 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=17425 $Y=18780 $D=1
M342 gnd! 265 249 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=17425 $Y=22270 $D=1
M343 gnd! 266 250 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=17425 $Y=25760 $D=1
M344 gnd! 267 251 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=17425 $Y=29250 $D=1
M345 gnd! 268 252 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=17425 $Y=32740 $D=1
M346 gnd! 269 253 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=17425 $Y=36230 $D=1
M347 gnd! 270 254 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=17425 $Y=39720 $D=1
M348 gnd! 271 255 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=17425 $Y=43210 $D=1
M349 gnd! 272 256 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=17425 $Y=46700 $D=1
M350 gnd! 273 257 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=17425 $Y=50190 $D=1
M351 gnd! 274 258 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=17425 $Y=53680 $D=1
M352 259 243 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=18015 $Y=1330 $D=1
M353 260 244 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=18015 $Y=4820 $D=1
M354 261 245 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=18015 $Y=8310 $D=1
M355 262 246 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=18015 $Y=11800 $D=1
M356 263 247 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=18015 $Y=15290 $D=1
M357 264 248 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=18015 $Y=18780 $D=1
M358 265 249 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=18015 $Y=22270 $D=1
M359 266 250 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=18015 $Y=25760 $D=1
M360 267 251 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=18015 $Y=29250 $D=1
M361 268 252 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=18015 $Y=32740 $D=1
M362 269 253 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=18015 $Y=36230 $D=1
M363 270 254 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=18015 $Y=39720 $D=1
M364 271 255 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=18015 $Y=43210 $D=1
M365 272 256 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=18015 $Y=46700 $D=1
M366 273 257 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=18015 $Y=50190 $D=1
M367 274 258 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=18015 $Y=53680 $D=1
M368 259 WL15 BL5 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=18455 $Y=1085 $D=1
M369 260 WL14 BL5 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=18455 $Y=4575 $D=1
M370 261 WL13 BL5 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=18455 $Y=8065 $D=1
M371 262 WL12 BL5 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=18455 $Y=11555 $D=1
M372 263 WL11 BL5 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=18455 $Y=15045 $D=1
M373 264 WL10 BL5 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=18455 $Y=18535 $D=1
M374 265 WL9 BL5 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=18455 $Y=22025 $D=1
M375 266 WL8 BL5 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=18455 $Y=25515 $D=1
M376 267 WL7 BL5 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=18455 $Y=29005 $D=1
M377 268 WL6 BL5 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=18455 $Y=32495 $D=1
M378 269 WL5 BL5 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=18455 $Y=35985 $D=1
M379 270 WL4 BL5 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=18455 $Y=39475 $D=1
M380 271 WL3 BL5 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=18455 $Y=42965 $D=1
M381 272 WL2 BL5 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=18455 $Y=46455 $D=1
M382 273 WL1 BL5 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=18455 $Y=49945 $D=1
M383 274 WL0 BL5 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=18455 $Y=53435 $D=1
M384 275 WL15 !BL6 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=19805 $Y=1085 $D=1
M385 276 WL14 !BL6 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=19805 $Y=4575 $D=1
M386 277 WL13 !BL6 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=19805 $Y=8065 $D=1
M387 278 WL12 !BL6 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=19805 $Y=11555 $D=1
M388 279 WL11 !BL6 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=19805 $Y=15045 $D=1
M389 280 WL10 !BL6 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=19805 $Y=18535 $D=1
M390 281 WL9 !BL6 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=19805 $Y=22025 $D=1
M391 282 WL8 !BL6 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=19805 $Y=25515 $D=1
M392 283 WL7 !BL6 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=19805 $Y=29005 $D=1
M393 284 WL6 !BL6 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=19805 $Y=32495 $D=1
M394 285 WL5 !BL6 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=19805 $Y=35985 $D=1
M395 286 WL4 !BL6 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=19805 $Y=39475 $D=1
M396 287 WL3 !BL6 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=19805 $Y=42965 $D=1
M397 288 WL2 !BL6 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=19805 $Y=46455 $D=1
M398 289 WL1 !BL6 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=19805 $Y=49945 $D=1
M399 290 WL0 !BL6 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=19805 $Y=53435 $D=1
M400 gnd! 291 275 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=20530 $Y=1330 $D=1
M401 gnd! 292 276 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=20530 $Y=4820 $D=1
M402 gnd! 293 277 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=20530 $Y=8310 $D=1
M403 gnd! 294 278 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=20530 $Y=11800 $D=1
M404 gnd! 295 279 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=20530 $Y=15290 $D=1
M405 gnd! 296 280 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=20530 $Y=18780 $D=1
M406 gnd! 297 281 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=20530 $Y=22270 $D=1
M407 gnd! 298 282 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=20530 $Y=25760 $D=1
M408 gnd! 299 283 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=20530 $Y=29250 $D=1
M409 gnd! 300 284 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=20530 $Y=32740 $D=1
M410 gnd! 301 285 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=20530 $Y=36230 $D=1
M411 gnd! 302 286 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=20530 $Y=39720 $D=1
M412 gnd! 303 287 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=20530 $Y=43210 $D=1
M413 gnd! 304 288 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=20530 $Y=46700 $D=1
M414 gnd! 305 289 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=20530 $Y=50190 $D=1
M415 gnd! 306 290 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=20530 $Y=53680 $D=1
M416 291 275 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=21120 $Y=1330 $D=1
M417 292 276 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=21120 $Y=4820 $D=1
M418 293 277 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=21120 $Y=8310 $D=1
M419 294 278 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=21120 $Y=11800 $D=1
M420 295 279 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=21120 $Y=15290 $D=1
M421 296 280 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=21120 $Y=18780 $D=1
M422 297 281 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=21120 $Y=22270 $D=1
M423 298 282 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=21120 $Y=25760 $D=1
M424 299 283 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=21120 $Y=29250 $D=1
M425 300 284 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=21120 $Y=32740 $D=1
M426 301 285 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=21120 $Y=36230 $D=1
M427 302 286 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=21120 $Y=39720 $D=1
M428 303 287 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=21120 $Y=43210 $D=1
M429 304 288 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=21120 $Y=46700 $D=1
M430 305 289 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=21120 $Y=50190 $D=1
M431 306 290 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=21120 $Y=53680 $D=1
M432 291 WL15 BL6 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=21560 $Y=1085 $D=1
M433 292 WL14 BL6 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=21560 $Y=4575 $D=1
M434 293 WL13 BL6 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=21560 $Y=8065 $D=1
M435 294 WL12 BL6 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=21560 $Y=11555 $D=1
M436 295 WL11 BL6 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=21560 $Y=15045 $D=1
M437 296 WL10 BL6 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=21560 $Y=18535 $D=1
M438 297 WL9 BL6 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=21560 $Y=22025 $D=1
M439 298 WL8 BL6 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=21560 $Y=25515 $D=1
M440 299 WL7 BL6 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=21560 $Y=29005 $D=1
M441 300 WL6 BL6 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=21560 $Y=32495 $D=1
M442 301 WL5 BL6 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=21560 $Y=35985 $D=1
M443 302 WL4 BL6 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=21560 $Y=39475 $D=1
M444 303 WL3 BL6 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=21560 $Y=42965 $D=1
M445 304 WL2 BL6 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=21560 $Y=46455 $D=1
M446 305 WL1 BL6 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=21560 $Y=49945 $D=1
M447 306 WL0 BL6 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=21560 $Y=53435 $D=1
M448 307 WL15 !BL7 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=22910 $Y=1085 $D=1
M449 308 WL14 !BL7 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=22910 $Y=4575 $D=1
M450 309 WL13 !BL7 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=22910 $Y=8065 $D=1
M451 310 WL12 !BL7 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=22910 $Y=11555 $D=1
M452 311 WL11 !BL7 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=22910 $Y=15045 $D=1
M453 312 WL10 !BL7 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=22910 $Y=18535 $D=1
M454 313 WL9 !BL7 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=22910 $Y=22025 $D=1
M455 314 WL8 !BL7 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=22910 $Y=25515 $D=1
M456 315 WL7 !BL7 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=22910 $Y=29005 $D=1
M457 316 WL6 !BL7 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=22910 $Y=32495 $D=1
M458 317 WL5 !BL7 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=22910 $Y=35985 $D=1
M459 318 WL4 !BL7 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=22910 $Y=39475 $D=1
M460 319 WL3 !BL7 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=22910 $Y=42965 $D=1
M461 320 WL2 !BL7 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=22910 $Y=46455 $D=1
M462 321 WL1 !BL7 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=22910 $Y=49945 $D=1
M463 322 WL0 !BL7 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=22910 $Y=53435 $D=1
M464 gnd! 323 307 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=23635 $Y=1330 $D=1
M465 gnd! 324 308 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=23635 $Y=4820 $D=1
M466 gnd! 325 309 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=23635 $Y=8310 $D=1
M467 gnd! 326 310 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=23635 $Y=11800 $D=1
M468 gnd! 327 311 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=23635 $Y=15290 $D=1
M469 gnd! 328 312 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=23635 $Y=18780 $D=1
M470 gnd! 329 313 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=23635 $Y=22270 $D=1
M471 gnd! 330 314 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=23635 $Y=25760 $D=1
M472 gnd! 331 315 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=23635 $Y=29250 $D=1
M473 gnd! 332 316 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=23635 $Y=32740 $D=1
M474 gnd! 333 317 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=23635 $Y=36230 $D=1
M475 gnd! 334 318 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=23635 $Y=39720 $D=1
M476 gnd! 335 319 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=23635 $Y=43210 $D=1
M477 gnd! 336 320 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=23635 $Y=46700 $D=1
M478 gnd! 337 321 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=23635 $Y=50190 $D=1
M479 gnd! 338 322 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=23635 $Y=53680 $D=1
M480 323 307 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=24225 $Y=1330 $D=1
M481 324 308 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=24225 $Y=4820 $D=1
M482 325 309 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=24225 $Y=8310 $D=1
M483 326 310 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=24225 $Y=11800 $D=1
M484 327 311 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=24225 $Y=15290 $D=1
M485 328 312 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=24225 $Y=18780 $D=1
M486 329 313 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=24225 $Y=22270 $D=1
M487 330 314 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=24225 $Y=25760 $D=1
M488 331 315 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=24225 $Y=29250 $D=1
M489 332 316 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=24225 $Y=32740 $D=1
M490 333 317 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=24225 $Y=36230 $D=1
M491 334 318 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=24225 $Y=39720 $D=1
M492 335 319 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=24225 $Y=43210 $D=1
M493 336 320 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=24225 $Y=46700 $D=1
M494 337 321 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=24225 $Y=50190 $D=1
M495 338 322 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=24225 $Y=53680 $D=1
M496 323 WL15 BL7 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=24665 $Y=1085 $D=1
M497 324 WL14 BL7 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=24665 $Y=4575 $D=1
M498 325 WL13 BL7 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=24665 $Y=8065 $D=1
M499 326 WL12 BL7 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=24665 $Y=11555 $D=1
M500 327 WL11 BL7 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=24665 $Y=15045 $D=1
M501 328 WL10 BL7 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=24665 $Y=18535 $D=1
M502 329 WL9 BL7 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=24665 $Y=22025 $D=1
M503 330 WL8 BL7 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=24665 $Y=25515 $D=1
M504 331 WL7 BL7 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=24665 $Y=29005 $D=1
M505 332 WL6 BL7 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=24665 $Y=32495 $D=1
M506 333 WL5 BL7 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=24665 $Y=35985 $D=1
M507 334 WL4 BL7 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=24665 $Y=39475 $D=1
M508 335 WL3 BL7 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=24665 $Y=42965 $D=1
M509 336 WL2 BL7 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=24665 $Y=46455 $D=1
M510 337 WL1 BL7 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=24665 $Y=49945 $D=1
M511 338 WL0 BL7 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=24665 $Y=53435 $D=1
M512 339 WL15 !BL8 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=26015 $Y=1085 $D=1
M513 340 WL14 !BL8 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=26015 $Y=4575 $D=1
M514 341 WL13 !BL8 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=26015 $Y=8065 $D=1
M515 342 WL12 !BL8 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=26015 $Y=11555 $D=1
M516 343 WL11 !BL8 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=26015 $Y=15045 $D=1
M517 344 WL10 !BL8 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=26015 $Y=18535 $D=1
M518 345 WL9 !BL8 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=26015 $Y=22025 $D=1
M519 346 WL8 !BL8 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=26015 $Y=25515 $D=1
M520 347 WL7 !BL8 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=26015 $Y=29005 $D=1
M521 348 WL6 !BL8 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=26015 $Y=32495 $D=1
M522 349 WL5 !BL8 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=26015 $Y=35985 $D=1
M523 350 WL4 !BL8 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=26015 $Y=39475 $D=1
M524 351 WL3 !BL8 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=26015 $Y=42965 $D=1
M525 352 WL2 !BL8 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=26015 $Y=46455 $D=1
M526 353 WL1 !BL8 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=26015 $Y=49945 $D=1
M527 354 WL0 !BL8 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=26015 $Y=53435 $D=1
M528 gnd! 355 339 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=26740 $Y=1330 $D=1
M529 gnd! 356 340 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=26740 $Y=4820 $D=1
M530 gnd! 357 341 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=26740 $Y=8310 $D=1
M531 gnd! 358 342 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=26740 $Y=11800 $D=1
M532 gnd! 359 343 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=26740 $Y=15290 $D=1
M533 gnd! 360 344 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=26740 $Y=18780 $D=1
M534 gnd! 361 345 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=26740 $Y=22270 $D=1
M535 gnd! 362 346 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=26740 $Y=25760 $D=1
M536 gnd! 363 347 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=26740 $Y=29250 $D=1
M537 gnd! 364 348 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=26740 $Y=32740 $D=1
M538 gnd! 365 349 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=26740 $Y=36230 $D=1
M539 gnd! 366 350 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=26740 $Y=39720 $D=1
M540 gnd! 367 351 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=26740 $Y=43210 $D=1
M541 gnd! 368 352 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=26740 $Y=46700 $D=1
M542 gnd! 369 353 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=26740 $Y=50190 $D=1
M543 gnd! 370 354 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=26740 $Y=53680 $D=1
M544 355 339 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=27330 $Y=1330 $D=1
M545 356 340 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=27330 $Y=4820 $D=1
M546 357 341 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=27330 $Y=8310 $D=1
M547 358 342 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=27330 $Y=11800 $D=1
M548 359 343 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=27330 $Y=15290 $D=1
M549 360 344 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=27330 $Y=18780 $D=1
M550 361 345 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=27330 $Y=22270 $D=1
M551 362 346 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=27330 $Y=25760 $D=1
M552 363 347 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=27330 $Y=29250 $D=1
M553 364 348 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=27330 $Y=32740 $D=1
M554 365 349 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=27330 $Y=36230 $D=1
M555 366 350 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=27330 $Y=39720 $D=1
M556 367 351 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=27330 $Y=43210 $D=1
M557 368 352 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=27330 $Y=46700 $D=1
M558 369 353 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=27330 $Y=50190 $D=1
M559 370 354 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=27330 $Y=53680 $D=1
M560 355 WL15 BL8 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=27770 $Y=1085 $D=1
M561 356 WL14 BL8 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=27770 $Y=4575 $D=1
M562 357 WL13 BL8 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=27770 $Y=8065 $D=1
M563 358 WL12 BL8 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=27770 $Y=11555 $D=1
M564 359 WL11 BL8 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=27770 $Y=15045 $D=1
M565 360 WL10 BL8 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=27770 $Y=18535 $D=1
M566 361 WL9 BL8 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=27770 $Y=22025 $D=1
M567 362 WL8 BL8 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=27770 $Y=25515 $D=1
M568 363 WL7 BL8 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=27770 $Y=29005 $D=1
M569 364 WL6 BL8 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=27770 $Y=32495 $D=1
M570 365 WL5 BL8 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=27770 $Y=35985 $D=1
M571 366 WL4 BL8 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=27770 $Y=39475 $D=1
M572 367 WL3 BL8 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=27770 $Y=42965 $D=1
M573 368 WL2 BL8 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=27770 $Y=46455 $D=1
M574 369 WL1 BL8 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=27770 $Y=49945 $D=1
M575 370 WL0 BL8 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=27770 $Y=53435 $D=1
M576 371 WL15 !BL9 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=29120 $Y=1085 $D=1
M577 372 WL14 !BL9 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=29120 $Y=4575 $D=1
M578 373 WL13 !BL9 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=29120 $Y=8065 $D=1
M579 374 WL12 !BL9 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=29120 $Y=11555 $D=1
M580 375 WL11 !BL9 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=29120 $Y=15045 $D=1
M581 376 WL10 !BL9 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=29120 $Y=18535 $D=1
M582 377 WL9 !BL9 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=29120 $Y=22025 $D=1
M583 378 WL8 !BL9 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=29120 $Y=25515 $D=1
M584 379 WL7 !BL9 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=29120 $Y=29005 $D=1
M585 380 WL6 !BL9 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=29120 $Y=32495 $D=1
M586 381 WL5 !BL9 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=29120 $Y=35985 $D=1
M587 382 WL4 !BL9 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=29120 $Y=39475 $D=1
M588 383 WL3 !BL9 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=29120 $Y=42965 $D=1
M589 384 WL2 !BL9 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=29120 $Y=46455 $D=1
M590 385 WL1 !BL9 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=29120 $Y=49945 $D=1
M591 386 WL0 !BL9 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=29120 $Y=53435 $D=1
M592 gnd! 387 371 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=29845 $Y=1330 $D=1
M593 gnd! 388 372 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=29845 $Y=4820 $D=1
M594 gnd! 389 373 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=29845 $Y=8310 $D=1
M595 gnd! 390 374 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=29845 $Y=11800 $D=1
M596 gnd! 391 375 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=29845 $Y=15290 $D=1
M597 gnd! 392 376 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=29845 $Y=18780 $D=1
M598 gnd! 393 377 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=29845 $Y=22270 $D=1
M599 gnd! 394 378 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=29845 $Y=25760 $D=1
M600 gnd! 395 379 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=29845 $Y=29250 $D=1
M601 gnd! 396 380 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=29845 $Y=32740 $D=1
M602 gnd! 397 381 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=29845 $Y=36230 $D=1
M603 gnd! 398 382 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=29845 $Y=39720 $D=1
M604 gnd! 399 383 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=29845 $Y=43210 $D=1
M605 gnd! 400 384 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=29845 $Y=46700 $D=1
M606 gnd! 401 385 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=29845 $Y=50190 $D=1
M607 gnd! 402 386 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=29845 $Y=53680 $D=1
M608 387 371 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=30435 $Y=1330 $D=1
M609 388 372 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=30435 $Y=4820 $D=1
M610 389 373 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=30435 $Y=8310 $D=1
M611 390 374 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=30435 $Y=11800 $D=1
M612 391 375 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=30435 $Y=15290 $D=1
M613 392 376 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=30435 $Y=18780 $D=1
M614 393 377 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=30435 $Y=22270 $D=1
M615 394 378 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=30435 $Y=25760 $D=1
M616 395 379 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=30435 $Y=29250 $D=1
M617 396 380 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=30435 $Y=32740 $D=1
M618 397 381 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=30435 $Y=36230 $D=1
M619 398 382 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=30435 $Y=39720 $D=1
M620 399 383 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=30435 $Y=43210 $D=1
M621 400 384 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=30435 $Y=46700 $D=1
M622 401 385 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=30435 $Y=50190 $D=1
M623 402 386 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=30435 $Y=53680 $D=1
M624 387 WL15 BL9 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=30875 $Y=1085 $D=1
M625 388 WL14 BL9 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=30875 $Y=4575 $D=1
M626 389 WL13 BL9 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=30875 $Y=8065 $D=1
M627 390 WL12 BL9 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=30875 $Y=11555 $D=1
M628 391 WL11 BL9 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=30875 $Y=15045 $D=1
M629 392 WL10 BL9 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=30875 $Y=18535 $D=1
M630 393 WL9 BL9 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=30875 $Y=22025 $D=1
M631 394 WL8 BL9 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=30875 $Y=25515 $D=1
M632 395 WL7 BL9 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=30875 $Y=29005 $D=1
M633 396 WL6 BL9 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=30875 $Y=32495 $D=1
M634 397 WL5 BL9 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=30875 $Y=35985 $D=1
M635 398 WL4 BL9 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=30875 $Y=39475 $D=1
M636 399 WL3 BL9 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=30875 $Y=42965 $D=1
M637 400 WL2 BL9 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=30875 $Y=46455 $D=1
M638 401 WL1 BL9 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=30875 $Y=49945 $D=1
M639 402 WL0 BL9 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=30875 $Y=53435 $D=1
M640 403 WL15 !BL10 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=32225 $Y=1085 $D=1
M641 404 WL14 !BL10 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=32225 $Y=4575 $D=1
M642 405 WL13 !BL10 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=32225 $Y=8065 $D=1
M643 406 WL12 !BL10 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=32225 $Y=11555 $D=1
M644 407 WL11 !BL10 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=32225 $Y=15045 $D=1
M645 408 WL10 !BL10 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=32225 $Y=18535 $D=1
M646 409 WL9 !BL10 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=32225 $Y=22025 $D=1
M647 410 WL8 !BL10 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=32225 $Y=25515 $D=1
M648 411 WL7 !BL10 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=32225 $Y=29005 $D=1
M649 412 WL6 !BL10 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=32225 $Y=32495 $D=1
M650 413 WL5 !BL10 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=32225 $Y=35985 $D=1
M651 414 WL4 !BL10 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=32225 $Y=39475 $D=1
M652 415 WL3 !BL10 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=32225 $Y=42965 $D=1
M653 416 WL2 !BL10 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=32225 $Y=46455 $D=1
M654 417 WL1 !BL10 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=32225 $Y=49945 $D=1
M655 418 WL0 !BL10 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=32225 $Y=53435 $D=1
M656 gnd! 419 403 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=32950 $Y=1330 $D=1
M657 gnd! 420 404 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=32950 $Y=4820 $D=1
M658 gnd! 421 405 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=32950 $Y=8310 $D=1
M659 gnd! 422 406 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=32950 $Y=11800 $D=1
M660 gnd! 423 407 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=32950 $Y=15290 $D=1
M661 gnd! 424 408 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=32950 $Y=18780 $D=1
M662 gnd! 425 409 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=32950 $Y=22270 $D=1
M663 gnd! 426 410 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=32950 $Y=25760 $D=1
M664 gnd! 427 411 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=32950 $Y=29250 $D=1
M665 gnd! 428 412 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=32950 $Y=32740 $D=1
M666 gnd! 429 413 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=32950 $Y=36230 $D=1
M667 gnd! 430 414 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=32950 $Y=39720 $D=1
M668 gnd! 431 415 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=32950 $Y=43210 $D=1
M669 gnd! 432 416 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=32950 $Y=46700 $D=1
M670 gnd! 433 417 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=32950 $Y=50190 $D=1
M671 gnd! 434 418 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=32950 $Y=53680 $D=1
M672 419 403 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=33540 $Y=1330 $D=1
M673 420 404 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=33540 $Y=4820 $D=1
M674 421 405 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=33540 $Y=8310 $D=1
M675 422 406 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=33540 $Y=11800 $D=1
M676 423 407 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=33540 $Y=15290 $D=1
M677 424 408 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=33540 $Y=18780 $D=1
M678 425 409 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=33540 $Y=22270 $D=1
M679 426 410 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=33540 $Y=25760 $D=1
M680 427 411 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=33540 $Y=29250 $D=1
M681 428 412 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=33540 $Y=32740 $D=1
M682 429 413 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=33540 $Y=36230 $D=1
M683 430 414 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=33540 $Y=39720 $D=1
M684 431 415 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=33540 $Y=43210 $D=1
M685 432 416 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=33540 $Y=46700 $D=1
M686 433 417 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=33540 $Y=50190 $D=1
M687 434 418 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=33540 $Y=53680 $D=1
M688 419 WL15 BL10 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=33980 $Y=1085 $D=1
M689 420 WL14 BL10 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=33980 $Y=4575 $D=1
M690 421 WL13 BL10 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=33980 $Y=8065 $D=1
M691 422 WL12 BL10 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=33980 $Y=11555 $D=1
M692 423 WL11 BL10 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=33980 $Y=15045 $D=1
M693 424 WL10 BL10 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=33980 $Y=18535 $D=1
M694 425 WL9 BL10 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=33980 $Y=22025 $D=1
M695 426 WL8 BL10 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=33980 $Y=25515 $D=1
M696 427 WL7 BL10 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=33980 $Y=29005 $D=1
M697 428 WL6 BL10 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=33980 $Y=32495 $D=1
M698 429 WL5 BL10 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=33980 $Y=35985 $D=1
M699 430 WL4 BL10 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=33980 $Y=39475 $D=1
M700 431 WL3 BL10 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=33980 $Y=42965 $D=1
M701 432 WL2 BL10 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=33980 $Y=46455 $D=1
M702 433 WL1 BL10 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=33980 $Y=49945 $D=1
M703 434 WL0 BL10 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=33980 $Y=53435 $D=1
M704 435 WL15 !BL11 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=35330 $Y=1085 $D=1
M705 436 WL14 !BL11 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=35330 $Y=4575 $D=1
M706 437 WL13 !BL11 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=35330 $Y=8065 $D=1
M707 438 WL12 !BL11 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=35330 $Y=11555 $D=1
M708 439 WL11 !BL11 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=35330 $Y=15045 $D=1
M709 440 WL10 !BL11 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=35330 $Y=18535 $D=1
M710 441 WL9 !BL11 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=35330 $Y=22025 $D=1
M711 442 WL8 !BL11 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=35330 $Y=25515 $D=1
M712 443 WL7 !BL11 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=35330 $Y=29005 $D=1
M713 444 WL6 !BL11 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=35330 $Y=32495 $D=1
M714 445 WL5 !BL11 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=35330 $Y=35985 $D=1
M715 446 WL4 !BL11 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=35330 $Y=39475 $D=1
M716 447 WL3 !BL11 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=35330 $Y=42965 $D=1
M717 448 WL2 !BL11 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=35330 $Y=46455 $D=1
M718 449 WL1 !BL11 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=35330 $Y=49945 $D=1
M719 450 WL0 !BL11 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=35330 $Y=53435 $D=1
M720 gnd! 451 435 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=36055 $Y=1330 $D=1
M721 gnd! 452 436 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=36055 $Y=4820 $D=1
M722 gnd! 453 437 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=36055 $Y=8310 $D=1
M723 gnd! 454 438 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=36055 $Y=11800 $D=1
M724 gnd! 455 439 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=36055 $Y=15290 $D=1
M725 gnd! 456 440 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=36055 $Y=18780 $D=1
M726 gnd! 457 441 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=36055 $Y=22270 $D=1
M727 gnd! 458 442 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=36055 $Y=25760 $D=1
M728 gnd! 459 443 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=36055 $Y=29250 $D=1
M729 gnd! 460 444 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=36055 $Y=32740 $D=1
M730 gnd! 461 445 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=36055 $Y=36230 $D=1
M731 gnd! 462 446 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=36055 $Y=39720 $D=1
M732 gnd! 463 447 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=36055 $Y=43210 $D=1
M733 gnd! 464 448 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=36055 $Y=46700 $D=1
M734 gnd! 465 449 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=36055 $Y=50190 $D=1
M735 gnd! 466 450 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=36055 $Y=53680 $D=1
M736 451 435 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=36645 $Y=1330 $D=1
M737 452 436 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=36645 $Y=4820 $D=1
M738 453 437 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=36645 $Y=8310 $D=1
M739 454 438 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=36645 $Y=11800 $D=1
M740 455 439 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=36645 $Y=15290 $D=1
M741 456 440 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=36645 $Y=18780 $D=1
M742 457 441 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=36645 $Y=22270 $D=1
M743 458 442 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=36645 $Y=25760 $D=1
M744 459 443 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=36645 $Y=29250 $D=1
M745 460 444 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=36645 $Y=32740 $D=1
M746 461 445 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=36645 $Y=36230 $D=1
M747 462 446 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=36645 $Y=39720 $D=1
M748 463 447 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=36645 $Y=43210 $D=1
M749 464 448 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=36645 $Y=46700 $D=1
M750 465 449 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=36645 $Y=50190 $D=1
M751 466 450 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=36645 $Y=53680 $D=1
M752 451 WL15 BL11 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=37085 $Y=1085 $D=1
M753 452 WL14 BL11 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=37085 $Y=4575 $D=1
M754 453 WL13 BL11 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=37085 $Y=8065 $D=1
M755 454 WL12 BL11 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=37085 $Y=11555 $D=1
M756 455 WL11 BL11 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=37085 $Y=15045 $D=1
M757 456 WL10 BL11 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=37085 $Y=18535 $D=1
M758 457 WL9 BL11 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=37085 $Y=22025 $D=1
M759 458 WL8 BL11 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=37085 $Y=25515 $D=1
M760 459 WL7 BL11 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=37085 $Y=29005 $D=1
M761 460 WL6 BL11 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=37085 $Y=32495 $D=1
M762 461 WL5 BL11 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=37085 $Y=35985 $D=1
M763 462 WL4 BL11 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=37085 $Y=39475 $D=1
M764 463 WL3 BL11 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=37085 $Y=42965 $D=1
M765 464 WL2 BL11 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=37085 $Y=46455 $D=1
M766 465 WL1 BL11 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=37085 $Y=49945 $D=1
M767 466 WL0 BL11 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=37085 $Y=53435 $D=1
M768 467 WL15 !BL12 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=38435 $Y=1085 $D=1
M769 468 WL14 !BL12 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=38435 $Y=4575 $D=1
M770 469 WL13 !BL12 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=38435 $Y=8065 $D=1
M771 470 WL12 !BL12 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=38435 $Y=11555 $D=1
M772 471 WL11 !BL12 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=38435 $Y=15045 $D=1
M773 472 WL10 !BL12 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=38435 $Y=18535 $D=1
M774 473 WL9 !BL12 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=38435 $Y=22025 $D=1
M775 474 WL8 !BL12 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=38435 $Y=25515 $D=1
M776 475 WL7 !BL12 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=38435 $Y=29005 $D=1
M777 476 WL6 !BL12 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=38435 $Y=32495 $D=1
M778 477 WL5 !BL12 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=38435 $Y=35985 $D=1
M779 478 WL4 !BL12 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=38435 $Y=39475 $D=1
M780 479 WL3 !BL12 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=38435 $Y=42965 $D=1
M781 480 WL2 !BL12 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=38435 $Y=46455 $D=1
M782 481 WL1 !BL12 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=38435 $Y=49945 $D=1
M783 482 WL0 !BL12 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=38435 $Y=53435 $D=1
M784 gnd! 483 467 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=39160 $Y=1330 $D=1
M785 gnd! 484 468 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=39160 $Y=4820 $D=1
M786 gnd! 485 469 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=39160 $Y=8310 $D=1
M787 gnd! 486 470 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=39160 $Y=11800 $D=1
M788 gnd! 487 471 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=39160 $Y=15290 $D=1
M789 gnd! 488 472 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=39160 $Y=18780 $D=1
M790 gnd! 489 473 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=39160 $Y=22270 $D=1
M791 gnd! 490 474 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=39160 $Y=25760 $D=1
M792 gnd! 491 475 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=39160 $Y=29250 $D=1
M793 gnd! 492 476 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=39160 $Y=32740 $D=1
M794 gnd! 493 477 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=39160 $Y=36230 $D=1
M795 gnd! 494 478 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=39160 $Y=39720 $D=1
M796 gnd! 495 479 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=39160 $Y=43210 $D=1
M797 gnd! 496 480 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=39160 $Y=46700 $D=1
M798 gnd! 497 481 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=39160 $Y=50190 $D=1
M799 gnd! 498 482 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=39160 $Y=53680 $D=1
M800 483 467 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=39750 $Y=1330 $D=1
M801 484 468 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=39750 $Y=4820 $D=1
M802 485 469 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=39750 $Y=8310 $D=1
M803 486 470 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=39750 $Y=11800 $D=1
M804 487 471 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=39750 $Y=15290 $D=1
M805 488 472 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=39750 $Y=18780 $D=1
M806 489 473 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=39750 $Y=22270 $D=1
M807 490 474 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=39750 $Y=25760 $D=1
M808 491 475 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=39750 $Y=29250 $D=1
M809 492 476 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=39750 $Y=32740 $D=1
M810 493 477 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=39750 $Y=36230 $D=1
M811 494 478 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=39750 $Y=39720 $D=1
M812 495 479 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=39750 $Y=43210 $D=1
M813 496 480 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=39750 $Y=46700 $D=1
M814 497 481 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=39750 $Y=50190 $D=1
M815 498 482 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=39750 $Y=53680 $D=1
M816 483 WL15 BL12 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=40190 $Y=1085 $D=1
M817 484 WL14 BL12 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=40190 $Y=4575 $D=1
M818 485 WL13 BL12 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=40190 $Y=8065 $D=1
M819 486 WL12 BL12 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=40190 $Y=11555 $D=1
M820 487 WL11 BL12 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=40190 $Y=15045 $D=1
M821 488 WL10 BL12 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=40190 $Y=18535 $D=1
M822 489 WL9 BL12 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=40190 $Y=22025 $D=1
M823 490 WL8 BL12 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=40190 $Y=25515 $D=1
M824 491 WL7 BL12 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=40190 $Y=29005 $D=1
M825 492 WL6 BL12 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=40190 $Y=32495 $D=1
M826 493 WL5 BL12 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=40190 $Y=35985 $D=1
M827 494 WL4 BL12 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=40190 $Y=39475 $D=1
M828 495 WL3 BL12 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=40190 $Y=42965 $D=1
M829 496 WL2 BL12 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=40190 $Y=46455 $D=1
M830 497 WL1 BL12 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=40190 $Y=49945 $D=1
M831 498 WL0 BL12 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=40190 $Y=53435 $D=1
M832 499 WL15 !BL13 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=41540 $Y=1085 $D=1
M833 500 WL14 !BL13 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=41540 $Y=4575 $D=1
M834 501 WL13 !BL13 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=41540 $Y=8065 $D=1
M835 502 WL12 !BL13 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=41540 $Y=11555 $D=1
M836 503 WL11 !BL13 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=41540 $Y=15045 $D=1
M837 504 WL10 !BL13 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=41540 $Y=18535 $D=1
M838 505 WL9 !BL13 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=41540 $Y=22025 $D=1
M839 506 WL8 !BL13 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=41540 $Y=25515 $D=1
M840 507 WL7 !BL13 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=41540 $Y=29005 $D=1
M841 508 WL6 !BL13 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=41540 $Y=32495 $D=1
M842 509 WL5 !BL13 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=41540 $Y=35985 $D=1
M843 510 WL4 !BL13 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=41540 $Y=39475 $D=1
M844 511 WL3 !BL13 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=41540 $Y=42965 $D=1
M845 512 WL2 !BL13 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=41540 $Y=46455 $D=1
M846 513 WL1 !BL13 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=41540 $Y=49945 $D=1
M847 514 WL0 !BL13 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=41540 $Y=53435 $D=1
M848 gnd! 515 499 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=42265 $Y=1330 $D=1
M849 gnd! 516 500 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=42265 $Y=4820 $D=1
M850 gnd! 517 501 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=42265 $Y=8310 $D=1
M851 gnd! 518 502 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=42265 $Y=11800 $D=1
M852 gnd! 519 503 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=42265 $Y=15290 $D=1
M853 gnd! 520 504 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=42265 $Y=18780 $D=1
M854 gnd! 521 505 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=42265 $Y=22270 $D=1
M855 gnd! 522 506 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=42265 $Y=25760 $D=1
M856 gnd! 523 507 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=42265 $Y=29250 $D=1
M857 gnd! 524 508 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=42265 $Y=32740 $D=1
M858 gnd! 525 509 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=42265 $Y=36230 $D=1
M859 gnd! 526 510 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=42265 $Y=39720 $D=1
M860 gnd! 527 511 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=42265 $Y=43210 $D=1
M861 gnd! 528 512 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=42265 $Y=46700 $D=1
M862 gnd! 529 513 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=42265 $Y=50190 $D=1
M863 gnd! 530 514 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=42265 $Y=53680 $D=1
M864 515 499 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=42855 $Y=1330 $D=1
M865 516 500 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=42855 $Y=4820 $D=1
M866 517 501 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=42855 $Y=8310 $D=1
M867 518 502 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=42855 $Y=11800 $D=1
M868 519 503 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=42855 $Y=15290 $D=1
M869 520 504 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=42855 $Y=18780 $D=1
M870 521 505 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=42855 $Y=22270 $D=1
M871 522 506 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=42855 $Y=25760 $D=1
M872 523 507 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=42855 $Y=29250 $D=1
M873 524 508 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=42855 $Y=32740 $D=1
M874 525 509 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=42855 $Y=36230 $D=1
M875 526 510 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=42855 $Y=39720 $D=1
M876 527 511 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=42855 $Y=43210 $D=1
M877 528 512 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=42855 $Y=46700 $D=1
M878 529 513 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=42855 $Y=50190 $D=1
M879 530 514 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=42855 $Y=53680 $D=1
M880 515 WL15 BL13 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=43295 $Y=1085 $D=1
M881 516 WL14 BL13 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=43295 $Y=4575 $D=1
M882 517 WL13 BL13 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=43295 $Y=8065 $D=1
M883 518 WL12 BL13 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=43295 $Y=11555 $D=1
M884 519 WL11 BL13 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=43295 $Y=15045 $D=1
M885 520 WL10 BL13 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=43295 $Y=18535 $D=1
M886 521 WL9 BL13 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=43295 $Y=22025 $D=1
M887 522 WL8 BL13 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=43295 $Y=25515 $D=1
M888 523 WL7 BL13 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=43295 $Y=29005 $D=1
M889 524 WL6 BL13 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=43295 $Y=32495 $D=1
M890 525 WL5 BL13 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=43295 $Y=35985 $D=1
M891 526 WL4 BL13 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=43295 $Y=39475 $D=1
M892 527 WL3 BL13 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=43295 $Y=42965 $D=1
M893 528 WL2 BL13 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=43295 $Y=46455 $D=1
M894 529 WL1 BL13 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=43295 $Y=49945 $D=1
M895 530 WL0 BL13 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=43295 $Y=53435 $D=1
M896 531 WL15 !BL14 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=44645 $Y=1085 $D=1
M897 532 WL14 !BL14 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=44645 $Y=4575 $D=1
M898 533 WL13 !BL14 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=44645 $Y=8065 $D=1
M899 534 WL12 !BL14 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=44645 $Y=11555 $D=1
M900 535 WL11 !BL14 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=44645 $Y=15045 $D=1
M901 536 WL10 !BL14 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=44645 $Y=18535 $D=1
M902 537 WL9 !BL14 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=44645 $Y=22025 $D=1
M903 538 WL8 !BL14 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=44645 $Y=25515 $D=1
M904 539 WL7 !BL14 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=44645 $Y=29005 $D=1
M905 540 WL6 !BL14 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=44645 $Y=32495 $D=1
M906 541 WL5 !BL14 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=44645 $Y=35985 $D=1
M907 542 WL4 !BL14 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=44645 $Y=39475 $D=1
M908 543 WL3 !BL14 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=44645 $Y=42965 $D=1
M909 544 WL2 !BL14 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=44645 $Y=46455 $D=1
M910 545 WL1 !BL14 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=44645 $Y=49945 $D=1
M911 546 WL0 !BL14 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=44645 $Y=53435 $D=1
M912 gnd! 547 531 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=45370 $Y=1330 $D=1
M913 gnd! 548 532 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=45370 $Y=4820 $D=1
M914 gnd! 549 533 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=45370 $Y=8310 $D=1
M915 gnd! 550 534 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=45370 $Y=11800 $D=1
M916 gnd! 551 535 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=45370 $Y=15290 $D=1
M917 gnd! 552 536 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=45370 $Y=18780 $D=1
M918 gnd! 553 537 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=45370 $Y=22270 $D=1
M919 gnd! 554 538 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=45370 $Y=25760 $D=1
M920 gnd! 555 539 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=45370 $Y=29250 $D=1
M921 gnd! 556 540 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=45370 $Y=32740 $D=1
M922 gnd! 557 541 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=45370 $Y=36230 $D=1
M923 gnd! 558 542 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=45370 $Y=39720 $D=1
M924 gnd! 559 543 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=45370 $Y=43210 $D=1
M925 gnd! 560 544 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=45370 $Y=46700 $D=1
M926 gnd! 561 545 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=45370 $Y=50190 $D=1
M927 gnd! 562 546 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=45370 $Y=53680 $D=1
M928 547 531 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=45960 $Y=1330 $D=1
M929 548 532 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=45960 $Y=4820 $D=1
M930 549 533 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=45960 $Y=8310 $D=1
M931 550 534 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=45960 $Y=11800 $D=1
M932 551 535 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=45960 $Y=15290 $D=1
M933 552 536 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=45960 $Y=18780 $D=1
M934 553 537 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=45960 $Y=22270 $D=1
M935 554 538 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=45960 $Y=25760 $D=1
M936 555 539 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=45960 $Y=29250 $D=1
M937 556 540 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=45960 $Y=32740 $D=1
M938 557 541 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=45960 $Y=36230 $D=1
M939 558 542 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=45960 $Y=39720 $D=1
M940 559 543 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=45960 $Y=43210 $D=1
M941 560 544 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=45960 $Y=46700 $D=1
M942 561 545 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=45960 $Y=50190 $D=1
M943 562 546 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=45960 $Y=53680 $D=1
M944 547 WL15 BL14 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=46400 $Y=1085 $D=1
M945 548 WL14 BL14 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=46400 $Y=4575 $D=1
M946 549 WL13 BL14 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=46400 $Y=8065 $D=1
M947 550 WL12 BL14 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=46400 $Y=11555 $D=1
M948 551 WL11 BL14 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=46400 $Y=15045 $D=1
M949 552 WL10 BL14 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=46400 $Y=18535 $D=1
M950 553 WL9 BL14 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=46400 $Y=22025 $D=1
M951 554 WL8 BL14 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=46400 $Y=25515 $D=1
M952 555 WL7 BL14 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=46400 $Y=29005 $D=1
M953 556 WL6 BL14 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=46400 $Y=32495 $D=1
M954 557 WL5 BL14 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=46400 $Y=35985 $D=1
M955 558 WL4 BL14 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=46400 $Y=39475 $D=1
M956 559 WL3 BL14 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=46400 $Y=42965 $D=1
M957 560 WL2 BL14 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=46400 $Y=46455 $D=1
M958 561 WL1 BL14 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=46400 $Y=49945 $D=1
M959 562 WL0 BL14 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=46400 $Y=53435 $D=1
M960 563 WL15 !BL15 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=47750 $Y=1085 $D=1
M961 564 WL14 !BL15 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=47750 $Y=4575 $D=1
M962 565 WL13 !BL15 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=47750 $Y=8065 $D=1
M963 566 WL12 !BL15 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=47750 $Y=11555 $D=1
M964 567 WL11 !BL15 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=47750 $Y=15045 $D=1
M965 568 WL10 !BL15 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=47750 $Y=18535 $D=1
M966 569 WL9 !BL15 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=47750 $Y=22025 $D=1
M967 570 WL8 !BL15 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=47750 $Y=25515 $D=1
M968 571 WL7 !BL15 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=47750 $Y=29005 $D=1
M969 572 WL6 !BL15 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=47750 $Y=32495 $D=1
M970 573 WL5 !BL15 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=47750 $Y=35985 $D=1
M971 574 WL4 !BL15 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=47750 $Y=39475 $D=1
M972 575 WL3 !BL15 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=47750 $Y=42965 $D=1
M973 576 WL2 !BL15 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=47750 $Y=46455 $D=1
M974 577 WL1 !BL15 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=47750 $Y=49945 $D=1
M975 578 WL0 !BL15 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=47750 $Y=53435 $D=1
M976 gnd! 579 563 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=48475 $Y=1330 $D=1
M977 gnd! 580 564 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=48475 $Y=4820 $D=1
M978 gnd! 581 565 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=48475 $Y=8310 $D=1
M979 gnd! 582 566 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=48475 $Y=11800 $D=1
M980 gnd! 583 567 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=48475 $Y=15290 $D=1
M981 gnd! 584 568 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=48475 $Y=18780 $D=1
M982 gnd! 585 569 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=48475 $Y=22270 $D=1
M983 gnd! 586 570 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=48475 $Y=25760 $D=1
M984 gnd! 587 571 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=48475 $Y=29250 $D=1
M985 gnd! 588 572 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=48475 $Y=32740 $D=1
M986 gnd! 589 573 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=48475 $Y=36230 $D=1
M987 gnd! 590 574 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=48475 $Y=39720 $D=1
M988 gnd! 591 575 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=48475 $Y=43210 $D=1
M989 gnd! 592 576 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=48475 $Y=46700 $D=1
M990 gnd! 593 577 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=48475 $Y=50190 $D=1
M991 gnd! 594 578 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=48475 $Y=53680 $D=1
M992 579 563 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=49065 $Y=1330 $D=1
M993 580 564 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=49065 $Y=4820 $D=1
M994 581 565 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=49065 $Y=8310 $D=1
M995 582 566 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=49065 $Y=11800 $D=1
M996 583 567 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=49065 $Y=15290 $D=1
M997 584 568 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=49065 $Y=18780 $D=1
M998 585 569 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=49065 $Y=22270 $D=1
M999 586 570 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=49065 $Y=25760 $D=1
M1000 587 571 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=49065 $Y=29250 $D=1
M1001 588 572 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=49065 $Y=32740 $D=1
M1002 589 573 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=49065 $Y=36230 $D=1
M1003 590 574 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=49065 $Y=39720 $D=1
M1004 591 575 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=49065 $Y=43210 $D=1
M1005 592 576 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=49065 $Y=46700 $D=1
M1006 593 577 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=49065 $Y=50190 $D=1
M1007 594 578 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=49065 $Y=53680 $D=1
M1008 579 WL15 BL15 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=49505 $Y=1085 $D=1
M1009 580 WL14 BL15 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=49505 $Y=4575 $D=1
M1010 581 WL13 BL15 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=49505 $Y=8065 $D=1
M1011 582 WL12 BL15 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=49505 $Y=11555 $D=1
M1012 583 WL11 BL15 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=49505 $Y=15045 $D=1
M1013 584 WL10 BL15 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=49505 $Y=18535 $D=1
M1014 585 WL9 BL15 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=49505 $Y=22025 $D=1
M1015 586 WL8 BL15 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=49505 $Y=25515 $D=1
M1016 587 WL7 BL15 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=49505 $Y=29005 $D=1
M1017 588 WL6 BL15 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=49505 $Y=32495 $D=1
M1018 589 WL5 BL15 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=49505 $Y=35985 $D=1
M1019 590 WL4 BL15 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=49505 $Y=39475 $D=1
M1020 591 WL3 BL15 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=49505 $Y=42965 $D=1
M1021 592 WL2 BL15 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=49505 $Y=46455 $D=1
M1022 593 WL1 BL15 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=49505 $Y=49945 $D=1
M1023 594 WL0 BL15 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=49505 $Y=53435 $D=1
M1024 595 WL15 !BL16 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=50855 $Y=1085 $D=1
M1025 596 WL14 !BL16 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=50855 $Y=4575 $D=1
M1026 597 WL13 !BL16 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=50855 $Y=8065 $D=1
M1027 598 WL12 !BL16 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=50855 $Y=11555 $D=1
M1028 599 WL11 !BL16 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=50855 $Y=15045 $D=1
M1029 600 WL10 !BL16 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=50855 $Y=18535 $D=1
M1030 601 WL9 !BL16 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=50855 $Y=22025 $D=1
M1031 602 WL8 !BL16 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=50855 $Y=25515 $D=1
M1032 603 WL7 !BL16 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=50855 $Y=29005 $D=1
M1033 604 WL6 !BL16 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=50855 $Y=32495 $D=1
M1034 605 WL5 !BL16 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=50855 $Y=35985 $D=1
M1035 606 WL4 !BL16 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=50855 $Y=39475 $D=1
M1036 607 WL3 !BL16 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=50855 $Y=42965 $D=1
M1037 608 WL2 !BL16 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=50855 $Y=46455 $D=1
M1038 609 WL1 !BL16 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=50855 $Y=49945 $D=1
M1039 610 WL0 !BL16 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=50855 $Y=53435 $D=1
M1040 gnd! 611 595 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=51580 $Y=1330 $D=1
M1041 gnd! 612 596 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=51580 $Y=4820 $D=1
M1042 gnd! 613 597 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=51580 $Y=8310 $D=1
M1043 gnd! 614 598 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=51580 $Y=11800 $D=1
M1044 gnd! 615 599 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=51580 $Y=15290 $D=1
M1045 gnd! 616 600 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=51580 $Y=18780 $D=1
M1046 gnd! 617 601 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=51580 $Y=22270 $D=1
M1047 gnd! 618 602 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=51580 $Y=25760 $D=1
M1048 gnd! 619 603 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=51580 $Y=29250 $D=1
M1049 gnd! 620 604 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=51580 $Y=32740 $D=1
M1050 gnd! 621 605 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=51580 $Y=36230 $D=1
M1051 gnd! 622 606 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=51580 $Y=39720 $D=1
M1052 gnd! 623 607 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=51580 $Y=43210 $D=1
M1053 gnd! 624 608 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=51580 $Y=46700 $D=1
M1054 gnd! 625 609 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=51580 $Y=50190 $D=1
M1055 gnd! 626 610 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=51580 $Y=53680 $D=1
M1056 611 595 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=52170 $Y=1330 $D=1
M1057 612 596 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=52170 $Y=4820 $D=1
M1058 613 597 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=52170 $Y=8310 $D=1
M1059 614 598 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=52170 $Y=11800 $D=1
M1060 615 599 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=52170 $Y=15290 $D=1
M1061 616 600 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=52170 $Y=18780 $D=1
M1062 617 601 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=52170 $Y=22270 $D=1
M1063 618 602 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=52170 $Y=25760 $D=1
M1064 619 603 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=52170 $Y=29250 $D=1
M1065 620 604 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=52170 $Y=32740 $D=1
M1066 621 605 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=52170 $Y=36230 $D=1
M1067 622 606 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=52170 $Y=39720 $D=1
M1068 623 607 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=52170 $Y=43210 $D=1
M1069 624 608 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=52170 $Y=46700 $D=1
M1070 625 609 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=52170 $Y=50190 $D=1
M1071 626 610 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=52170 $Y=53680 $D=1
M1072 611 WL15 BL16 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=52610 $Y=1085 $D=1
M1073 612 WL14 BL16 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=52610 $Y=4575 $D=1
M1074 613 WL13 BL16 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=52610 $Y=8065 $D=1
M1075 614 WL12 BL16 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=52610 $Y=11555 $D=1
M1076 615 WL11 BL16 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=52610 $Y=15045 $D=1
M1077 616 WL10 BL16 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=52610 $Y=18535 $D=1
M1078 617 WL9 BL16 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=52610 $Y=22025 $D=1
M1079 618 WL8 BL16 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=52610 $Y=25515 $D=1
M1080 619 WL7 BL16 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=52610 $Y=29005 $D=1
M1081 620 WL6 BL16 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=52610 $Y=32495 $D=1
M1082 621 WL5 BL16 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=52610 $Y=35985 $D=1
M1083 622 WL4 BL16 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=52610 $Y=39475 $D=1
M1084 623 WL3 BL16 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=52610 $Y=42965 $D=1
M1085 624 WL2 BL16 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=52610 $Y=46455 $D=1
M1086 625 WL1 BL16 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=52610 $Y=49945 $D=1
M1087 626 WL0 BL16 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=52610 $Y=53435 $D=1
M1088 627 WL15 !BL17 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=53960 $Y=1085 $D=1
M1089 628 WL14 !BL17 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=53960 $Y=4575 $D=1
M1090 629 WL13 !BL17 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=53960 $Y=8065 $D=1
M1091 630 WL12 !BL17 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=53960 $Y=11555 $D=1
M1092 631 WL11 !BL17 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=53960 $Y=15045 $D=1
M1093 632 WL10 !BL17 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=53960 $Y=18535 $D=1
M1094 633 WL9 !BL17 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=53960 $Y=22025 $D=1
M1095 634 WL8 !BL17 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=53960 $Y=25515 $D=1
M1096 635 WL7 !BL17 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=53960 $Y=29005 $D=1
M1097 636 WL6 !BL17 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=53960 $Y=32495 $D=1
M1098 637 WL5 !BL17 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=53960 $Y=35985 $D=1
M1099 638 WL4 !BL17 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=53960 $Y=39475 $D=1
M1100 639 WL3 !BL17 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=53960 $Y=42965 $D=1
M1101 640 WL2 !BL17 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=53960 $Y=46455 $D=1
M1102 641 WL1 !BL17 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=53960 $Y=49945 $D=1
M1103 642 WL0 !BL17 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=53960 $Y=53435 $D=1
M1104 gnd! 643 627 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=54685 $Y=1330 $D=1
M1105 gnd! 644 628 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=54685 $Y=4820 $D=1
M1106 gnd! 645 629 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=54685 $Y=8310 $D=1
M1107 gnd! 646 630 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=54685 $Y=11800 $D=1
M1108 gnd! 647 631 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=54685 $Y=15290 $D=1
M1109 gnd! 648 632 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=54685 $Y=18780 $D=1
M1110 gnd! 649 633 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=54685 $Y=22270 $D=1
M1111 gnd! 650 634 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=54685 $Y=25760 $D=1
M1112 gnd! 651 635 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=54685 $Y=29250 $D=1
M1113 gnd! 652 636 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=54685 $Y=32740 $D=1
M1114 gnd! 653 637 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=54685 $Y=36230 $D=1
M1115 gnd! 654 638 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=54685 $Y=39720 $D=1
M1116 gnd! 655 639 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=54685 $Y=43210 $D=1
M1117 gnd! 656 640 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=54685 $Y=46700 $D=1
M1118 gnd! 657 641 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=54685 $Y=50190 $D=1
M1119 gnd! 658 642 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=54685 $Y=53680 $D=1
M1120 643 627 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=55275 $Y=1330 $D=1
M1121 644 628 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=55275 $Y=4820 $D=1
M1122 645 629 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=55275 $Y=8310 $D=1
M1123 646 630 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=55275 $Y=11800 $D=1
M1124 647 631 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=55275 $Y=15290 $D=1
M1125 648 632 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=55275 $Y=18780 $D=1
M1126 649 633 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=55275 $Y=22270 $D=1
M1127 650 634 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=55275 $Y=25760 $D=1
M1128 651 635 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=55275 $Y=29250 $D=1
M1129 652 636 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=55275 $Y=32740 $D=1
M1130 653 637 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=55275 $Y=36230 $D=1
M1131 654 638 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=55275 $Y=39720 $D=1
M1132 655 639 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=55275 $Y=43210 $D=1
M1133 656 640 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=55275 $Y=46700 $D=1
M1134 657 641 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=55275 $Y=50190 $D=1
M1135 658 642 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=55275 $Y=53680 $D=1
M1136 643 WL15 BL17 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=55715 $Y=1085 $D=1
M1137 644 WL14 BL17 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=55715 $Y=4575 $D=1
M1138 645 WL13 BL17 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=55715 $Y=8065 $D=1
M1139 646 WL12 BL17 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=55715 $Y=11555 $D=1
M1140 647 WL11 BL17 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=55715 $Y=15045 $D=1
M1141 648 WL10 BL17 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=55715 $Y=18535 $D=1
M1142 649 WL9 BL17 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=55715 $Y=22025 $D=1
M1143 650 WL8 BL17 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=55715 $Y=25515 $D=1
M1144 651 WL7 BL17 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=55715 $Y=29005 $D=1
M1145 652 WL6 BL17 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=55715 $Y=32495 $D=1
M1146 653 WL5 BL17 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=55715 $Y=35985 $D=1
M1147 654 WL4 BL17 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=55715 $Y=39475 $D=1
M1148 655 WL3 BL17 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=55715 $Y=42965 $D=1
M1149 656 WL2 BL17 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=55715 $Y=46455 $D=1
M1150 657 WL1 BL17 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=55715 $Y=49945 $D=1
M1151 658 WL0 BL17 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=55715 $Y=53435 $D=1
M1152 659 WL15 !BL18 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=57065 $Y=1085 $D=1
M1153 660 WL14 !BL18 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=57065 $Y=4575 $D=1
M1154 661 WL13 !BL18 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=57065 $Y=8065 $D=1
M1155 662 WL12 !BL18 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=57065 $Y=11555 $D=1
M1156 663 WL11 !BL18 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=57065 $Y=15045 $D=1
M1157 664 WL10 !BL18 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=57065 $Y=18535 $D=1
M1158 665 WL9 !BL18 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=57065 $Y=22025 $D=1
M1159 666 WL8 !BL18 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=57065 $Y=25515 $D=1
M1160 667 WL7 !BL18 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=57065 $Y=29005 $D=1
M1161 668 WL6 !BL18 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=57065 $Y=32495 $D=1
M1162 669 WL5 !BL18 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=57065 $Y=35985 $D=1
M1163 670 WL4 !BL18 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=57065 $Y=39475 $D=1
M1164 671 WL3 !BL18 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=57065 $Y=42965 $D=1
M1165 672 WL2 !BL18 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=57065 $Y=46455 $D=1
M1166 673 WL1 !BL18 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=57065 $Y=49945 $D=1
M1167 674 WL0 !BL18 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=57065 $Y=53435 $D=1
M1168 gnd! 675 659 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=57790 $Y=1330 $D=1
M1169 gnd! 676 660 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=57790 $Y=4820 $D=1
M1170 gnd! 677 661 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=57790 $Y=8310 $D=1
M1171 gnd! 678 662 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=57790 $Y=11800 $D=1
M1172 gnd! 679 663 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=57790 $Y=15290 $D=1
M1173 gnd! 680 664 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=57790 $Y=18780 $D=1
M1174 gnd! 681 665 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=57790 $Y=22270 $D=1
M1175 gnd! 682 666 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=57790 $Y=25760 $D=1
M1176 gnd! 683 667 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=57790 $Y=29250 $D=1
M1177 gnd! 684 668 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=57790 $Y=32740 $D=1
M1178 gnd! 685 669 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=57790 $Y=36230 $D=1
M1179 gnd! 686 670 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=57790 $Y=39720 $D=1
M1180 gnd! 687 671 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=57790 $Y=43210 $D=1
M1181 gnd! 688 672 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=57790 $Y=46700 $D=1
M1182 gnd! 689 673 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=57790 $Y=50190 $D=1
M1183 gnd! 690 674 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=57790 $Y=53680 $D=1
M1184 675 659 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=58380 $Y=1330 $D=1
M1185 676 660 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=58380 $Y=4820 $D=1
M1186 677 661 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=58380 $Y=8310 $D=1
M1187 678 662 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=58380 $Y=11800 $D=1
M1188 679 663 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=58380 $Y=15290 $D=1
M1189 680 664 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=58380 $Y=18780 $D=1
M1190 681 665 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=58380 $Y=22270 $D=1
M1191 682 666 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=58380 $Y=25760 $D=1
M1192 683 667 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=58380 $Y=29250 $D=1
M1193 684 668 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=58380 $Y=32740 $D=1
M1194 685 669 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=58380 $Y=36230 $D=1
M1195 686 670 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=58380 $Y=39720 $D=1
M1196 687 671 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=58380 $Y=43210 $D=1
M1197 688 672 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=58380 $Y=46700 $D=1
M1198 689 673 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=58380 $Y=50190 $D=1
M1199 690 674 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=58380 $Y=53680 $D=1
M1200 675 WL15 BL18 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=58820 $Y=1085 $D=1
M1201 676 WL14 BL18 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=58820 $Y=4575 $D=1
M1202 677 WL13 BL18 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=58820 $Y=8065 $D=1
M1203 678 WL12 BL18 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=58820 $Y=11555 $D=1
M1204 679 WL11 BL18 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=58820 $Y=15045 $D=1
M1205 680 WL10 BL18 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=58820 $Y=18535 $D=1
M1206 681 WL9 BL18 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=58820 $Y=22025 $D=1
M1207 682 WL8 BL18 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=58820 $Y=25515 $D=1
M1208 683 WL7 BL18 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=58820 $Y=29005 $D=1
M1209 684 WL6 BL18 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=58820 $Y=32495 $D=1
M1210 685 WL5 BL18 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=58820 $Y=35985 $D=1
M1211 686 WL4 BL18 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=58820 $Y=39475 $D=1
M1212 687 WL3 BL18 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=58820 $Y=42965 $D=1
M1213 688 WL2 BL18 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=58820 $Y=46455 $D=1
M1214 689 WL1 BL18 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=58820 $Y=49945 $D=1
M1215 690 WL0 BL18 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=58820 $Y=53435 $D=1
M1216 691 WL15 !BL19 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=60170 $Y=1085 $D=1
M1217 692 WL14 !BL19 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=60170 $Y=4575 $D=1
M1218 693 WL13 !BL19 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=60170 $Y=8065 $D=1
M1219 694 WL12 !BL19 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=60170 $Y=11555 $D=1
M1220 695 WL11 !BL19 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=60170 $Y=15045 $D=1
M1221 696 WL10 !BL19 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=60170 $Y=18535 $D=1
M1222 697 WL9 !BL19 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=60170 $Y=22025 $D=1
M1223 698 WL8 !BL19 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=60170 $Y=25515 $D=1
M1224 699 WL7 !BL19 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=60170 $Y=29005 $D=1
M1225 700 WL6 !BL19 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=60170 $Y=32495 $D=1
M1226 701 WL5 !BL19 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=60170 $Y=35985 $D=1
M1227 702 WL4 !BL19 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=60170 $Y=39475 $D=1
M1228 703 WL3 !BL19 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=60170 $Y=42965 $D=1
M1229 704 WL2 !BL19 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=60170 $Y=46455 $D=1
M1230 705 WL1 !BL19 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=60170 $Y=49945 $D=1
M1231 706 WL0 !BL19 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=60170 $Y=53435 $D=1
M1232 gnd! 707 691 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=60895 $Y=1330 $D=1
M1233 gnd! 708 692 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=60895 $Y=4820 $D=1
M1234 gnd! 709 693 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=60895 $Y=8310 $D=1
M1235 gnd! 710 694 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=60895 $Y=11800 $D=1
M1236 gnd! 711 695 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=60895 $Y=15290 $D=1
M1237 gnd! 712 696 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=60895 $Y=18780 $D=1
M1238 gnd! 713 697 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=60895 $Y=22270 $D=1
M1239 gnd! 714 698 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=60895 $Y=25760 $D=1
M1240 gnd! 715 699 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=60895 $Y=29250 $D=1
M1241 gnd! 716 700 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=60895 $Y=32740 $D=1
M1242 gnd! 717 701 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=60895 $Y=36230 $D=1
M1243 gnd! 718 702 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=60895 $Y=39720 $D=1
M1244 gnd! 719 703 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=60895 $Y=43210 $D=1
M1245 gnd! 720 704 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=60895 $Y=46700 $D=1
M1246 gnd! 721 705 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=60895 $Y=50190 $D=1
M1247 gnd! 722 706 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=60895 $Y=53680 $D=1
M1248 707 691 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=61485 $Y=1330 $D=1
M1249 708 692 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=61485 $Y=4820 $D=1
M1250 709 693 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=61485 $Y=8310 $D=1
M1251 710 694 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=61485 $Y=11800 $D=1
M1252 711 695 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=61485 $Y=15290 $D=1
M1253 712 696 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=61485 $Y=18780 $D=1
M1254 713 697 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=61485 $Y=22270 $D=1
M1255 714 698 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=61485 $Y=25760 $D=1
M1256 715 699 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=61485 $Y=29250 $D=1
M1257 716 700 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=61485 $Y=32740 $D=1
M1258 717 701 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=61485 $Y=36230 $D=1
M1259 718 702 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=61485 $Y=39720 $D=1
M1260 719 703 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=61485 $Y=43210 $D=1
M1261 720 704 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=61485 $Y=46700 $D=1
M1262 721 705 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=61485 $Y=50190 $D=1
M1263 722 706 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=61485 $Y=53680 $D=1
M1264 707 WL15 BL19 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=61925 $Y=1085 $D=1
M1265 708 WL14 BL19 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=61925 $Y=4575 $D=1
M1266 709 WL13 BL19 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=61925 $Y=8065 $D=1
M1267 710 WL12 BL19 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=61925 $Y=11555 $D=1
M1268 711 WL11 BL19 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=61925 $Y=15045 $D=1
M1269 712 WL10 BL19 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=61925 $Y=18535 $D=1
M1270 713 WL9 BL19 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=61925 $Y=22025 $D=1
M1271 714 WL8 BL19 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=61925 $Y=25515 $D=1
M1272 715 WL7 BL19 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=61925 $Y=29005 $D=1
M1273 716 WL6 BL19 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=61925 $Y=32495 $D=1
M1274 717 WL5 BL19 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=61925 $Y=35985 $D=1
M1275 718 WL4 BL19 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=61925 $Y=39475 $D=1
M1276 719 WL3 BL19 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=61925 $Y=42965 $D=1
M1277 720 WL2 BL19 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=61925 $Y=46455 $D=1
M1278 721 WL1 BL19 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=61925 $Y=49945 $D=1
M1279 722 WL0 BL19 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=61925 $Y=53435 $D=1
M1280 723 WL15 !BL20 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=63275 $Y=1085 $D=1
M1281 724 WL14 !BL20 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=63275 $Y=4575 $D=1
M1282 725 WL13 !BL20 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=63275 $Y=8065 $D=1
M1283 726 WL12 !BL20 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=63275 $Y=11555 $D=1
M1284 727 WL11 !BL20 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=63275 $Y=15045 $D=1
M1285 728 WL10 !BL20 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=63275 $Y=18535 $D=1
M1286 729 WL9 !BL20 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=63275 $Y=22025 $D=1
M1287 730 WL8 !BL20 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=63275 $Y=25515 $D=1
M1288 731 WL7 !BL20 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=63275 $Y=29005 $D=1
M1289 732 WL6 !BL20 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=63275 $Y=32495 $D=1
M1290 733 WL5 !BL20 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=63275 $Y=35985 $D=1
M1291 734 WL4 !BL20 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=63275 $Y=39475 $D=1
M1292 735 WL3 !BL20 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=63275 $Y=42965 $D=1
M1293 736 WL2 !BL20 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=63275 $Y=46455 $D=1
M1294 737 WL1 !BL20 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=63275 $Y=49945 $D=1
M1295 738 WL0 !BL20 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=63275 $Y=53435 $D=1
M1296 gnd! 739 723 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=64000 $Y=1330 $D=1
M1297 gnd! 740 724 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=64000 $Y=4820 $D=1
M1298 gnd! 741 725 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=64000 $Y=8310 $D=1
M1299 gnd! 742 726 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=64000 $Y=11800 $D=1
M1300 gnd! 743 727 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=64000 $Y=15290 $D=1
M1301 gnd! 744 728 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=64000 $Y=18780 $D=1
M1302 gnd! 745 729 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=64000 $Y=22270 $D=1
M1303 gnd! 746 730 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=64000 $Y=25760 $D=1
M1304 gnd! 747 731 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=64000 $Y=29250 $D=1
M1305 gnd! 748 732 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=64000 $Y=32740 $D=1
M1306 gnd! 749 733 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=64000 $Y=36230 $D=1
M1307 gnd! 750 734 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=64000 $Y=39720 $D=1
M1308 gnd! 751 735 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=64000 $Y=43210 $D=1
M1309 gnd! 752 736 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=64000 $Y=46700 $D=1
M1310 gnd! 753 737 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=64000 $Y=50190 $D=1
M1311 gnd! 754 738 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=64000 $Y=53680 $D=1
M1312 739 723 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=64590 $Y=1330 $D=1
M1313 740 724 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=64590 $Y=4820 $D=1
M1314 741 725 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=64590 $Y=8310 $D=1
M1315 742 726 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=64590 $Y=11800 $D=1
M1316 743 727 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=64590 $Y=15290 $D=1
M1317 744 728 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=64590 $Y=18780 $D=1
M1318 745 729 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=64590 $Y=22270 $D=1
M1319 746 730 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=64590 $Y=25760 $D=1
M1320 747 731 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=64590 $Y=29250 $D=1
M1321 748 732 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=64590 $Y=32740 $D=1
M1322 749 733 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=64590 $Y=36230 $D=1
M1323 750 734 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=64590 $Y=39720 $D=1
M1324 751 735 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=64590 $Y=43210 $D=1
M1325 752 736 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=64590 $Y=46700 $D=1
M1326 753 737 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=64590 $Y=50190 $D=1
M1327 754 738 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=64590 $Y=53680 $D=1
M1328 739 WL15 BL20 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=65030 $Y=1085 $D=1
M1329 740 WL14 BL20 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=65030 $Y=4575 $D=1
M1330 741 WL13 BL20 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=65030 $Y=8065 $D=1
M1331 742 WL12 BL20 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=65030 $Y=11555 $D=1
M1332 743 WL11 BL20 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=65030 $Y=15045 $D=1
M1333 744 WL10 BL20 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=65030 $Y=18535 $D=1
M1334 745 WL9 BL20 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=65030 $Y=22025 $D=1
M1335 746 WL8 BL20 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=65030 $Y=25515 $D=1
M1336 747 WL7 BL20 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=65030 $Y=29005 $D=1
M1337 748 WL6 BL20 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=65030 $Y=32495 $D=1
M1338 749 WL5 BL20 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=65030 $Y=35985 $D=1
M1339 750 WL4 BL20 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=65030 $Y=39475 $D=1
M1340 751 WL3 BL20 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=65030 $Y=42965 $D=1
M1341 752 WL2 BL20 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=65030 $Y=46455 $D=1
M1342 753 WL1 BL20 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=65030 $Y=49945 $D=1
M1343 754 WL0 BL20 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=65030 $Y=53435 $D=1
M1344 755 WL15 !BL21 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=66380 $Y=1085 $D=1
M1345 756 WL14 !BL21 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=66380 $Y=4575 $D=1
M1346 757 WL13 !BL21 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=66380 $Y=8065 $D=1
M1347 758 WL12 !BL21 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=66380 $Y=11555 $D=1
M1348 759 WL11 !BL21 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=66380 $Y=15045 $D=1
M1349 760 WL10 !BL21 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=66380 $Y=18535 $D=1
M1350 761 WL9 !BL21 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=66380 $Y=22025 $D=1
M1351 762 WL8 !BL21 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=66380 $Y=25515 $D=1
M1352 763 WL7 !BL21 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=66380 $Y=29005 $D=1
M1353 764 WL6 !BL21 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=66380 $Y=32495 $D=1
M1354 765 WL5 !BL21 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=66380 $Y=35985 $D=1
M1355 766 WL4 !BL21 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=66380 $Y=39475 $D=1
M1356 767 WL3 !BL21 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=66380 $Y=42965 $D=1
M1357 768 WL2 !BL21 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=66380 $Y=46455 $D=1
M1358 769 WL1 !BL21 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=66380 $Y=49945 $D=1
M1359 770 WL0 !BL21 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=66380 $Y=53435 $D=1
M1360 gnd! 771 755 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=67105 $Y=1330 $D=1
M1361 gnd! 772 756 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=67105 $Y=4820 $D=1
M1362 gnd! 773 757 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=67105 $Y=8310 $D=1
M1363 gnd! 774 758 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=67105 $Y=11800 $D=1
M1364 gnd! 775 759 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=67105 $Y=15290 $D=1
M1365 gnd! 776 760 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=67105 $Y=18780 $D=1
M1366 gnd! 777 761 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=67105 $Y=22270 $D=1
M1367 gnd! 778 762 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=67105 $Y=25760 $D=1
M1368 gnd! 779 763 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=67105 $Y=29250 $D=1
M1369 gnd! 780 764 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=67105 $Y=32740 $D=1
M1370 gnd! 781 765 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=67105 $Y=36230 $D=1
M1371 gnd! 782 766 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=67105 $Y=39720 $D=1
M1372 gnd! 783 767 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=67105 $Y=43210 $D=1
M1373 gnd! 784 768 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=67105 $Y=46700 $D=1
M1374 gnd! 785 769 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=67105 $Y=50190 $D=1
M1375 gnd! 786 770 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=67105 $Y=53680 $D=1
M1376 771 755 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=67695 $Y=1330 $D=1
M1377 772 756 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=67695 $Y=4820 $D=1
M1378 773 757 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=67695 $Y=8310 $D=1
M1379 774 758 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=67695 $Y=11800 $D=1
M1380 775 759 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=67695 $Y=15290 $D=1
M1381 776 760 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=67695 $Y=18780 $D=1
M1382 777 761 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=67695 $Y=22270 $D=1
M1383 778 762 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=67695 $Y=25760 $D=1
M1384 779 763 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=67695 $Y=29250 $D=1
M1385 780 764 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=67695 $Y=32740 $D=1
M1386 781 765 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=67695 $Y=36230 $D=1
M1387 782 766 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=67695 $Y=39720 $D=1
M1388 783 767 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=67695 $Y=43210 $D=1
M1389 784 768 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=67695 $Y=46700 $D=1
M1390 785 769 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=67695 $Y=50190 $D=1
M1391 786 770 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=67695 $Y=53680 $D=1
M1392 771 WL15 BL21 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=68135 $Y=1085 $D=1
M1393 772 WL14 BL21 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=68135 $Y=4575 $D=1
M1394 773 WL13 BL21 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=68135 $Y=8065 $D=1
M1395 774 WL12 BL21 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=68135 $Y=11555 $D=1
M1396 775 WL11 BL21 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=68135 $Y=15045 $D=1
M1397 776 WL10 BL21 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=68135 $Y=18535 $D=1
M1398 777 WL9 BL21 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=68135 $Y=22025 $D=1
M1399 778 WL8 BL21 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=68135 $Y=25515 $D=1
M1400 779 WL7 BL21 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=68135 $Y=29005 $D=1
M1401 780 WL6 BL21 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=68135 $Y=32495 $D=1
M1402 781 WL5 BL21 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=68135 $Y=35985 $D=1
M1403 782 WL4 BL21 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=68135 $Y=39475 $D=1
M1404 783 WL3 BL21 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=68135 $Y=42965 $D=1
M1405 784 WL2 BL21 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=68135 $Y=46455 $D=1
M1406 785 WL1 BL21 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=68135 $Y=49945 $D=1
M1407 786 WL0 BL21 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=68135 $Y=53435 $D=1
M1408 787 WL15 !BL22 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=69485 $Y=1085 $D=1
M1409 788 WL14 !BL22 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=69485 $Y=4575 $D=1
M1410 789 WL13 !BL22 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=69485 $Y=8065 $D=1
M1411 790 WL12 !BL22 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=69485 $Y=11555 $D=1
M1412 791 WL11 !BL22 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=69485 $Y=15045 $D=1
M1413 792 WL10 !BL22 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=69485 $Y=18535 $D=1
M1414 793 WL9 !BL22 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=69485 $Y=22025 $D=1
M1415 794 WL8 !BL22 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=69485 $Y=25515 $D=1
M1416 795 WL7 !BL22 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=69485 $Y=29005 $D=1
M1417 796 WL6 !BL22 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=69485 $Y=32495 $D=1
M1418 797 WL5 !BL22 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=69485 $Y=35985 $D=1
M1419 798 WL4 !BL22 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=69485 $Y=39475 $D=1
M1420 799 WL3 !BL22 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=69485 $Y=42965 $D=1
M1421 800 WL2 !BL22 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=69485 $Y=46455 $D=1
M1422 801 WL1 !BL22 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=69485 $Y=49945 $D=1
M1423 802 WL0 !BL22 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=69485 $Y=53435 $D=1
M1424 gnd! 803 787 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=70210 $Y=1330 $D=1
M1425 gnd! 804 788 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=70210 $Y=4820 $D=1
M1426 gnd! 805 789 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=70210 $Y=8310 $D=1
M1427 gnd! 806 790 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=70210 $Y=11800 $D=1
M1428 gnd! 807 791 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=70210 $Y=15290 $D=1
M1429 gnd! 808 792 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=70210 $Y=18780 $D=1
M1430 gnd! 809 793 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=70210 $Y=22270 $D=1
M1431 gnd! 810 794 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=70210 $Y=25760 $D=1
M1432 gnd! 811 795 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=70210 $Y=29250 $D=1
M1433 gnd! 812 796 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=70210 $Y=32740 $D=1
M1434 gnd! 813 797 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=70210 $Y=36230 $D=1
M1435 gnd! 814 798 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=70210 $Y=39720 $D=1
M1436 gnd! 815 799 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=70210 $Y=43210 $D=1
M1437 gnd! 816 800 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=70210 $Y=46700 $D=1
M1438 gnd! 817 801 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=70210 $Y=50190 $D=1
M1439 gnd! 818 802 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=70210 $Y=53680 $D=1
M1440 803 787 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=70800 $Y=1330 $D=1
M1441 804 788 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=70800 $Y=4820 $D=1
M1442 805 789 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=70800 $Y=8310 $D=1
M1443 806 790 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=70800 $Y=11800 $D=1
M1444 807 791 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=70800 $Y=15290 $D=1
M1445 808 792 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=70800 $Y=18780 $D=1
M1446 809 793 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=70800 $Y=22270 $D=1
M1447 810 794 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=70800 $Y=25760 $D=1
M1448 811 795 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=70800 $Y=29250 $D=1
M1449 812 796 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=70800 $Y=32740 $D=1
M1450 813 797 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=70800 $Y=36230 $D=1
M1451 814 798 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=70800 $Y=39720 $D=1
M1452 815 799 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=70800 $Y=43210 $D=1
M1453 816 800 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=70800 $Y=46700 $D=1
M1454 817 801 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=70800 $Y=50190 $D=1
M1455 818 802 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=70800 $Y=53680 $D=1
M1456 803 WL15 BL22 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=71240 $Y=1085 $D=1
M1457 804 WL14 BL22 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=71240 $Y=4575 $D=1
M1458 805 WL13 BL22 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=71240 $Y=8065 $D=1
M1459 806 WL12 BL22 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=71240 $Y=11555 $D=1
M1460 807 WL11 BL22 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=71240 $Y=15045 $D=1
M1461 808 WL10 BL22 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=71240 $Y=18535 $D=1
M1462 809 WL9 BL22 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=71240 $Y=22025 $D=1
M1463 810 WL8 BL22 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=71240 $Y=25515 $D=1
M1464 811 WL7 BL22 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=71240 $Y=29005 $D=1
M1465 812 WL6 BL22 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=71240 $Y=32495 $D=1
M1466 813 WL5 BL22 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=71240 $Y=35985 $D=1
M1467 814 WL4 BL22 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=71240 $Y=39475 $D=1
M1468 815 WL3 BL22 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=71240 $Y=42965 $D=1
M1469 816 WL2 BL22 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=71240 $Y=46455 $D=1
M1470 817 WL1 BL22 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=71240 $Y=49945 $D=1
M1471 818 WL0 BL22 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=71240 $Y=53435 $D=1
M1472 819 WL15 !BL23 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=72590 $Y=1085 $D=1
M1473 820 WL14 !BL23 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=72590 $Y=4575 $D=1
M1474 821 WL13 !BL23 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=72590 $Y=8065 $D=1
M1475 822 WL12 !BL23 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=72590 $Y=11555 $D=1
M1476 823 WL11 !BL23 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=72590 $Y=15045 $D=1
M1477 824 WL10 !BL23 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=72590 $Y=18535 $D=1
M1478 825 WL9 !BL23 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=72590 $Y=22025 $D=1
M1479 826 WL8 !BL23 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=72590 $Y=25515 $D=1
M1480 827 WL7 !BL23 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=72590 $Y=29005 $D=1
M1481 828 WL6 !BL23 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=72590 $Y=32495 $D=1
M1482 829 WL5 !BL23 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=72590 $Y=35985 $D=1
M1483 830 WL4 !BL23 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=72590 $Y=39475 $D=1
M1484 831 WL3 !BL23 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=72590 $Y=42965 $D=1
M1485 832 WL2 !BL23 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=72590 $Y=46455 $D=1
M1486 833 WL1 !BL23 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=72590 $Y=49945 $D=1
M1487 834 WL0 !BL23 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=72590 $Y=53435 $D=1
M1488 gnd! 835 819 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=73315 $Y=1330 $D=1
M1489 gnd! 836 820 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=73315 $Y=4820 $D=1
M1490 gnd! 837 821 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=73315 $Y=8310 $D=1
M1491 gnd! 838 822 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=73315 $Y=11800 $D=1
M1492 gnd! 839 823 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=73315 $Y=15290 $D=1
M1493 gnd! 840 824 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=73315 $Y=18780 $D=1
M1494 gnd! 841 825 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=73315 $Y=22270 $D=1
M1495 gnd! 842 826 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=73315 $Y=25760 $D=1
M1496 gnd! 843 827 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=73315 $Y=29250 $D=1
M1497 gnd! 844 828 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=73315 $Y=32740 $D=1
M1498 gnd! 845 829 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=73315 $Y=36230 $D=1
M1499 gnd! 846 830 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=73315 $Y=39720 $D=1
M1500 gnd! 847 831 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=73315 $Y=43210 $D=1
M1501 gnd! 848 832 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=73315 $Y=46700 $D=1
M1502 gnd! 849 833 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=73315 $Y=50190 $D=1
M1503 gnd! 850 834 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=73315 $Y=53680 $D=1
M1504 835 819 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=73905 $Y=1330 $D=1
M1505 836 820 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=73905 $Y=4820 $D=1
M1506 837 821 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=73905 $Y=8310 $D=1
M1507 838 822 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=73905 $Y=11800 $D=1
M1508 839 823 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=73905 $Y=15290 $D=1
M1509 840 824 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=73905 $Y=18780 $D=1
M1510 841 825 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=73905 $Y=22270 $D=1
M1511 842 826 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=73905 $Y=25760 $D=1
M1512 843 827 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=73905 $Y=29250 $D=1
M1513 844 828 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=73905 $Y=32740 $D=1
M1514 845 829 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=73905 $Y=36230 $D=1
M1515 846 830 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=73905 $Y=39720 $D=1
M1516 847 831 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=73905 $Y=43210 $D=1
M1517 848 832 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=73905 $Y=46700 $D=1
M1518 849 833 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=73905 $Y=50190 $D=1
M1519 850 834 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=73905 $Y=53680 $D=1
M1520 835 WL15 BL23 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=74345 $Y=1085 $D=1
M1521 836 WL14 BL23 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=74345 $Y=4575 $D=1
M1522 837 WL13 BL23 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=74345 $Y=8065 $D=1
M1523 838 WL12 BL23 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=74345 $Y=11555 $D=1
M1524 839 WL11 BL23 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=74345 $Y=15045 $D=1
M1525 840 WL10 BL23 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=74345 $Y=18535 $D=1
M1526 841 WL9 BL23 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=74345 $Y=22025 $D=1
M1527 842 WL8 BL23 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=74345 $Y=25515 $D=1
M1528 843 WL7 BL23 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=74345 $Y=29005 $D=1
M1529 844 WL6 BL23 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=74345 $Y=32495 $D=1
M1530 845 WL5 BL23 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=74345 $Y=35985 $D=1
M1531 846 WL4 BL23 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=74345 $Y=39475 $D=1
M1532 847 WL3 BL23 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=74345 $Y=42965 $D=1
M1533 848 WL2 BL23 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=74345 $Y=46455 $D=1
M1534 849 WL1 BL23 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=74345 $Y=49945 $D=1
M1535 850 WL0 BL23 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=74345 $Y=53435 $D=1
M1536 851 WL15 !BL24 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=75695 $Y=1085 $D=1
M1537 852 WL14 !BL24 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=75695 $Y=4575 $D=1
M1538 853 WL13 !BL24 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=75695 $Y=8065 $D=1
M1539 854 WL12 !BL24 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=75695 $Y=11555 $D=1
M1540 855 WL11 !BL24 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=75695 $Y=15045 $D=1
M1541 856 WL10 !BL24 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=75695 $Y=18535 $D=1
M1542 857 WL9 !BL24 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=75695 $Y=22025 $D=1
M1543 858 WL8 !BL24 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=75695 $Y=25515 $D=1
M1544 859 WL7 !BL24 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=75695 $Y=29005 $D=1
M1545 860 WL6 !BL24 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=75695 $Y=32495 $D=1
M1546 861 WL5 !BL24 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=75695 $Y=35985 $D=1
M1547 862 WL4 !BL24 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=75695 $Y=39475 $D=1
M1548 863 WL3 !BL24 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=75695 $Y=42965 $D=1
M1549 864 WL2 !BL24 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=75695 $Y=46455 $D=1
M1550 865 WL1 !BL24 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=75695 $Y=49945 $D=1
M1551 866 WL0 !BL24 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=75695 $Y=53435 $D=1
M1552 gnd! 867 851 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=76420 $Y=1330 $D=1
M1553 gnd! 868 852 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=76420 $Y=4820 $D=1
M1554 gnd! 869 853 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=76420 $Y=8310 $D=1
M1555 gnd! 870 854 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=76420 $Y=11800 $D=1
M1556 gnd! 871 855 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=76420 $Y=15290 $D=1
M1557 gnd! 872 856 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=76420 $Y=18780 $D=1
M1558 gnd! 873 857 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=76420 $Y=22270 $D=1
M1559 gnd! 874 858 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=76420 $Y=25760 $D=1
M1560 gnd! 875 859 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=76420 $Y=29250 $D=1
M1561 gnd! 876 860 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=76420 $Y=32740 $D=1
M1562 gnd! 877 861 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=76420 $Y=36230 $D=1
M1563 gnd! 878 862 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=76420 $Y=39720 $D=1
M1564 gnd! 879 863 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=76420 $Y=43210 $D=1
M1565 gnd! 880 864 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=76420 $Y=46700 $D=1
M1566 gnd! 881 865 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=76420 $Y=50190 $D=1
M1567 gnd! 882 866 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=76420 $Y=53680 $D=1
M1568 867 851 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=77010 $Y=1330 $D=1
M1569 868 852 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=77010 $Y=4820 $D=1
M1570 869 853 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=77010 $Y=8310 $D=1
M1571 870 854 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=77010 $Y=11800 $D=1
M1572 871 855 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=77010 $Y=15290 $D=1
M1573 872 856 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=77010 $Y=18780 $D=1
M1574 873 857 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=77010 $Y=22270 $D=1
M1575 874 858 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=77010 $Y=25760 $D=1
M1576 875 859 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=77010 $Y=29250 $D=1
M1577 876 860 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=77010 $Y=32740 $D=1
M1578 877 861 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=77010 $Y=36230 $D=1
M1579 878 862 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=77010 $Y=39720 $D=1
M1580 879 863 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=77010 $Y=43210 $D=1
M1581 880 864 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=77010 $Y=46700 $D=1
M1582 881 865 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=77010 $Y=50190 $D=1
M1583 882 866 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=77010 $Y=53680 $D=1
M1584 867 WL15 BL24 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=77450 $Y=1085 $D=1
M1585 868 WL14 BL24 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=77450 $Y=4575 $D=1
M1586 869 WL13 BL24 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=77450 $Y=8065 $D=1
M1587 870 WL12 BL24 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=77450 $Y=11555 $D=1
M1588 871 WL11 BL24 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=77450 $Y=15045 $D=1
M1589 872 WL10 BL24 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=77450 $Y=18535 $D=1
M1590 873 WL9 BL24 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=77450 $Y=22025 $D=1
M1591 874 WL8 BL24 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=77450 $Y=25515 $D=1
M1592 875 WL7 BL24 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=77450 $Y=29005 $D=1
M1593 876 WL6 BL24 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=77450 $Y=32495 $D=1
M1594 877 WL5 BL24 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=77450 $Y=35985 $D=1
M1595 878 WL4 BL24 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=77450 $Y=39475 $D=1
M1596 879 WL3 BL24 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=77450 $Y=42965 $D=1
M1597 880 WL2 BL24 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=77450 $Y=46455 $D=1
M1598 881 WL1 BL24 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=77450 $Y=49945 $D=1
M1599 882 WL0 BL24 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=77450 $Y=53435 $D=1
M1600 883 WL15 !BL25 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=78800 $Y=1085 $D=1
M1601 884 WL14 !BL25 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=78800 $Y=4575 $D=1
M1602 885 WL13 !BL25 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=78800 $Y=8065 $D=1
M1603 886 WL12 !BL25 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=78800 $Y=11555 $D=1
M1604 887 WL11 !BL25 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=78800 $Y=15045 $D=1
M1605 888 WL10 !BL25 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=78800 $Y=18535 $D=1
M1606 889 WL9 !BL25 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=78800 $Y=22025 $D=1
M1607 890 WL8 !BL25 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=78800 $Y=25515 $D=1
M1608 891 WL7 !BL25 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=78800 $Y=29005 $D=1
M1609 892 WL6 !BL25 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=78800 $Y=32495 $D=1
M1610 893 WL5 !BL25 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=78800 $Y=35985 $D=1
M1611 894 WL4 !BL25 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=78800 $Y=39475 $D=1
M1612 895 WL3 !BL25 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=78800 $Y=42965 $D=1
M1613 896 WL2 !BL25 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=78800 $Y=46455 $D=1
M1614 897 WL1 !BL25 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=78800 $Y=49945 $D=1
M1615 898 WL0 !BL25 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=78800 $Y=53435 $D=1
M1616 gnd! 899 883 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=79525 $Y=1330 $D=1
M1617 gnd! 900 884 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=79525 $Y=4820 $D=1
M1618 gnd! 901 885 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=79525 $Y=8310 $D=1
M1619 gnd! 902 886 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=79525 $Y=11800 $D=1
M1620 gnd! 903 887 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=79525 $Y=15290 $D=1
M1621 gnd! 904 888 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=79525 $Y=18780 $D=1
M1622 gnd! 905 889 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=79525 $Y=22270 $D=1
M1623 gnd! 906 890 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=79525 $Y=25760 $D=1
M1624 gnd! 907 891 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=79525 $Y=29250 $D=1
M1625 gnd! 908 892 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=79525 $Y=32740 $D=1
M1626 gnd! 909 893 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=79525 $Y=36230 $D=1
M1627 gnd! 910 894 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=79525 $Y=39720 $D=1
M1628 gnd! 911 895 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=79525 $Y=43210 $D=1
M1629 gnd! 912 896 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=79525 $Y=46700 $D=1
M1630 gnd! 913 897 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=79525 $Y=50190 $D=1
M1631 gnd! 914 898 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=79525 $Y=53680 $D=1
M1632 899 883 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=80115 $Y=1330 $D=1
M1633 900 884 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=80115 $Y=4820 $D=1
M1634 901 885 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=80115 $Y=8310 $D=1
M1635 902 886 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=80115 $Y=11800 $D=1
M1636 903 887 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=80115 $Y=15290 $D=1
M1637 904 888 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=80115 $Y=18780 $D=1
M1638 905 889 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=80115 $Y=22270 $D=1
M1639 906 890 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=80115 $Y=25760 $D=1
M1640 907 891 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=80115 $Y=29250 $D=1
M1641 908 892 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=80115 $Y=32740 $D=1
M1642 909 893 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=80115 $Y=36230 $D=1
M1643 910 894 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=80115 $Y=39720 $D=1
M1644 911 895 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=80115 $Y=43210 $D=1
M1645 912 896 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=80115 $Y=46700 $D=1
M1646 913 897 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=80115 $Y=50190 $D=1
M1647 914 898 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=80115 $Y=53680 $D=1
M1648 899 WL15 BL25 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=80555 $Y=1085 $D=1
M1649 900 WL14 BL25 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=80555 $Y=4575 $D=1
M1650 901 WL13 BL25 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=80555 $Y=8065 $D=1
M1651 902 WL12 BL25 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=80555 $Y=11555 $D=1
M1652 903 WL11 BL25 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=80555 $Y=15045 $D=1
M1653 904 WL10 BL25 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=80555 $Y=18535 $D=1
M1654 905 WL9 BL25 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=80555 $Y=22025 $D=1
M1655 906 WL8 BL25 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=80555 $Y=25515 $D=1
M1656 907 WL7 BL25 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=80555 $Y=29005 $D=1
M1657 908 WL6 BL25 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=80555 $Y=32495 $D=1
M1658 909 WL5 BL25 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=80555 $Y=35985 $D=1
M1659 910 WL4 BL25 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=80555 $Y=39475 $D=1
M1660 911 WL3 BL25 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=80555 $Y=42965 $D=1
M1661 912 WL2 BL25 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=80555 $Y=46455 $D=1
M1662 913 WL1 BL25 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=80555 $Y=49945 $D=1
M1663 914 WL0 BL25 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=80555 $Y=53435 $D=1
M1664 915 WL15 !BL26 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=81905 $Y=1085 $D=1
M1665 916 WL14 !BL26 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=81905 $Y=4575 $D=1
M1666 917 WL13 !BL26 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=81905 $Y=8065 $D=1
M1667 918 WL12 !BL26 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=81905 $Y=11555 $D=1
M1668 919 WL11 !BL26 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=81905 $Y=15045 $D=1
M1669 920 WL10 !BL26 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=81905 $Y=18535 $D=1
M1670 921 WL9 !BL26 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=81905 $Y=22025 $D=1
M1671 922 WL8 !BL26 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=81905 $Y=25515 $D=1
M1672 923 WL7 !BL26 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=81905 $Y=29005 $D=1
M1673 924 WL6 !BL26 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=81905 $Y=32495 $D=1
M1674 925 WL5 !BL26 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=81905 $Y=35985 $D=1
M1675 926 WL4 !BL26 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=81905 $Y=39475 $D=1
M1676 927 WL3 !BL26 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=81905 $Y=42965 $D=1
M1677 928 WL2 !BL26 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=81905 $Y=46455 $D=1
M1678 929 WL1 !BL26 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=81905 $Y=49945 $D=1
M1679 930 WL0 !BL26 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=81905 $Y=53435 $D=1
M1680 gnd! 931 915 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=82630 $Y=1330 $D=1
M1681 gnd! 932 916 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=82630 $Y=4820 $D=1
M1682 gnd! 933 917 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=82630 $Y=8310 $D=1
M1683 gnd! 934 918 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=82630 $Y=11800 $D=1
M1684 gnd! 935 919 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=82630 $Y=15290 $D=1
M1685 gnd! 936 920 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=82630 $Y=18780 $D=1
M1686 gnd! 937 921 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=82630 $Y=22270 $D=1
M1687 gnd! 938 922 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=82630 $Y=25760 $D=1
M1688 gnd! 939 923 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=82630 $Y=29250 $D=1
M1689 gnd! 940 924 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=82630 $Y=32740 $D=1
M1690 gnd! 941 925 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=82630 $Y=36230 $D=1
M1691 gnd! 942 926 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=82630 $Y=39720 $D=1
M1692 gnd! 943 927 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=82630 $Y=43210 $D=1
M1693 gnd! 944 928 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=82630 $Y=46700 $D=1
M1694 gnd! 945 929 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=82630 $Y=50190 $D=1
M1695 gnd! 946 930 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=82630 $Y=53680 $D=1
M1696 931 915 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=83220 $Y=1330 $D=1
M1697 932 916 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=83220 $Y=4820 $D=1
M1698 933 917 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=83220 $Y=8310 $D=1
M1699 934 918 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=83220 $Y=11800 $D=1
M1700 935 919 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=83220 $Y=15290 $D=1
M1701 936 920 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=83220 $Y=18780 $D=1
M1702 937 921 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=83220 $Y=22270 $D=1
M1703 938 922 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=83220 $Y=25760 $D=1
M1704 939 923 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=83220 $Y=29250 $D=1
M1705 940 924 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=83220 $Y=32740 $D=1
M1706 941 925 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=83220 $Y=36230 $D=1
M1707 942 926 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=83220 $Y=39720 $D=1
M1708 943 927 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=83220 $Y=43210 $D=1
M1709 944 928 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=83220 $Y=46700 $D=1
M1710 945 929 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=83220 $Y=50190 $D=1
M1711 946 930 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=83220 $Y=53680 $D=1
M1712 931 WL15 BL26 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=83660 $Y=1085 $D=1
M1713 932 WL14 BL26 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=83660 $Y=4575 $D=1
M1714 933 WL13 BL26 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=83660 $Y=8065 $D=1
M1715 934 WL12 BL26 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=83660 $Y=11555 $D=1
M1716 935 WL11 BL26 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=83660 $Y=15045 $D=1
M1717 936 WL10 BL26 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=83660 $Y=18535 $D=1
M1718 937 WL9 BL26 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=83660 $Y=22025 $D=1
M1719 938 WL8 BL26 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=83660 $Y=25515 $D=1
M1720 939 WL7 BL26 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=83660 $Y=29005 $D=1
M1721 940 WL6 BL26 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=83660 $Y=32495 $D=1
M1722 941 WL5 BL26 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=83660 $Y=35985 $D=1
M1723 942 WL4 BL26 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=83660 $Y=39475 $D=1
M1724 943 WL3 BL26 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=83660 $Y=42965 $D=1
M1725 944 WL2 BL26 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=83660 $Y=46455 $D=1
M1726 945 WL1 BL26 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=83660 $Y=49945 $D=1
M1727 946 WL0 BL26 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=83660 $Y=53435 $D=1
M1728 947 WL15 !BL27 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=85010 $Y=1085 $D=1
M1729 948 WL14 !BL27 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=85010 $Y=4575 $D=1
M1730 949 WL13 !BL27 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=85010 $Y=8065 $D=1
M1731 950 WL12 !BL27 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=85010 $Y=11555 $D=1
M1732 951 WL11 !BL27 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=85010 $Y=15045 $D=1
M1733 952 WL10 !BL27 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=85010 $Y=18535 $D=1
M1734 953 WL9 !BL27 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=85010 $Y=22025 $D=1
M1735 954 WL8 !BL27 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=85010 $Y=25515 $D=1
M1736 955 WL7 !BL27 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=85010 $Y=29005 $D=1
M1737 956 WL6 !BL27 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=85010 $Y=32495 $D=1
M1738 957 WL5 !BL27 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=85010 $Y=35985 $D=1
M1739 958 WL4 !BL27 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=85010 $Y=39475 $D=1
M1740 959 WL3 !BL27 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=85010 $Y=42965 $D=1
M1741 960 WL2 !BL27 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=85010 $Y=46455 $D=1
M1742 961 WL1 !BL27 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=85010 $Y=49945 $D=1
M1743 962 WL0 !BL27 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=85010 $Y=53435 $D=1
M1744 gnd! 963 947 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=85735 $Y=1330 $D=1
M1745 gnd! 964 948 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=85735 $Y=4820 $D=1
M1746 gnd! 965 949 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=85735 $Y=8310 $D=1
M1747 gnd! 966 950 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=85735 $Y=11800 $D=1
M1748 gnd! 967 951 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=85735 $Y=15290 $D=1
M1749 gnd! 968 952 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=85735 $Y=18780 $D=1
M1750 gnd! 969 953 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=85735 $Y=22270 $D=1
M1751 gnd! 970 954 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=85735 $Y=25760 $D=1
M1752 gnd! 971 955 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=85735 $Y=29250 $D=1
M1753 gnd! 972 956 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=85735 $Y=32740 $D=1
M1754 gnd! 973 957 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=85735 $Y=36230 $D=1
M1755 gnd! 974 958 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=85735 $Y=39720 $D=1
M1756 gnd! 975 959 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=85735 $Y=43210 $D=1
M1757 gnd! 976 960 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=85735 $Y=46700 $D=1
M1758 gnd! 977 961 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=85735 $Y=50190 $D=1
M1759 gnd! 978 962 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=85735 $Y=53680 $D=1
M1760 963 947 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=86325 $Y=1330 $D=1
M1761 964 948 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=86325 $Y=4820 $D=1
M1762 965 949 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=86325 $Y=8310 $D=1
M1763 966 950 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=86325 $Y=11800 $D=1
M1764 967 951 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=86325 $Y=15290 $D=1
M1765 968 952 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=86325 $Y=18780 $D=1
M1766 969 953 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=86325 $Y=22270 $D=1
M1767 970 954 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=86325 $Y=25760 $D=1
M1768 971 955 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=86325 $Y=29250 $D=1
M1769 972 956 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=86325 $Y=32740 $D=1
M1770 973 957 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=86325 $Y=36230 $D=1
M1771 974 958 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=86325 $Y=39720 $D=1
M1772 975 959 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=86325 $Y=43210 $D=1
M1773 976 960 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=86325 $Y=46700 $D=1
M1774 977 961 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=86325 $Y=50190 $D=1
M1775 978 962 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=86325 $Y=53680 $D=1
M1776 963 WL15 BL27 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=86765 $Y=1085 $D=1
M1777 964 WL14 BL27 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=86765 $Y=4575 $D=1
M1778 965 WL13 BL27 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=86765 $Y=8065 $D=1
M1779 966 WL12 BL27 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=86765 $Y=11555 $D=1
M1780 967 WL11 BL27 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=86765 $Y=15045 $D=1
M1781 968 WL10 BL27 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=86765 $Y=18535 $D=1
M1782 969 WL9 BL27 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=86765 $Y=22025 $D=1
M1783 970 WL8 BL27 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=86765 $Y=25515 $D=1
M1784 971 WL7 BL27 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=86765 $Y=29005 $D=1
M1785 972 WL6 BL27 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=86765 $Y=32495 $D=1
M1786 973 WL5 BL27 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=86765 $Y=35985 $D=1
M1787 974 WL4 BL27 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=86765 $Y=39475 $D=1
M1788 975 WL3 BL27 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=86765 $Y=42965 $D=1
M1789 976 WL2 BL27 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=86765 $Y=46455 $D=1
M1790 977 WL1 BL27 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=86765 $Y=49945 $D=1
M1791 978 WL0 BL27 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=86765 $Y=53435 $D=1
M1792 979 WL15 !BL28 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=88115 $Y=1085 $D=1
M1793 980 WL14 !BL28 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=88115 $Y=4575 $D=1
M1794 981 WL13 !BL28 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=88115 $Y=8065 $D=1
M1795 982 WL12 !BL28 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=88115 $Y=11555 $D=1
M1796 983 WL11 !BL28 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=88115 $Y=15045 $D=1
M1797 984 WL10 !BL28 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=88115 $Y=18535 $D=1
M1798 985 WL9 !BL28 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=88115 $Y=22025 $D=1
M1799 986 WL8 !BL28 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=88115 $Y=25515 $D=1
M1800 987 WL7 !BL28 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=88115 $Y=29005 $D=1
M1801 988 WL6 !BL28 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=88115 $Y=32495 $D=1
M1802 989 WL5 !BL28 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=88115 $Y=35985 $D=1
M1803 990 WL4 !BL28 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=88115 $Y=39475 $D=1
M1804 991 WL3 !BL28 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=88115 $Y=42965 $D=1
M1805 992 WL2 !BL28 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=88115 $Y=46455 $D=1
M1806 993 WL1 !BL28 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=88115 $Y=49945 $D=1
M1807 994 WL0 !BL28 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=88115 $Y=53435 $D=1
M1808 gnd! 995 979 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=88840 $Y=1330 $D=1
M1809 gnd! 996 980 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=88840 $Y=4820 $D=1
M1810 gnd! 997 981 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=88840 $Y=8310 $D=1
M1811 gnd! 998 982 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=88840 $Y=11800 $D=1
M1812 gnd! 999 983 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=88840 $Y=15290 $D=1
M1813 gnd! 1000 984 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=88840 $Y=18780 $D=1
M1814 gnd! 1001 985 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=88840 $Y=22270 $D=1
M1815 gnd! 1002 986 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=88840 $Y=25760 $D=1
M1816 gnd! 1003 987 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=88840 $Y=29250 $D=1
M1817 gnd! 1004 988 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=88840 $Y=32740 $D=1
M1818 gnd! 1005 989 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=88840 $Y=36230 $D=1
M1819 gnd! 1006 990 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=88840 $Y=39720 $D=1
M1820 gnd! 1007 991 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=88840 $Y=43210 $D=1
M1821 gnd! 1008 992 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=88840 $Y=46700 $D=1
M1822 gnd! 1009 993 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=88840 $Y=50190 $D=1
M1823 gnd! 1010 994 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=88840 $Y=53680 $D=1
M1824 995 979 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=89430 $Y=1330 $D=1
M1825 996 980 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=89430 $Y=4820 $D=1
M1826 997 981 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=89430 $Y=8310 $D=1
M1827 998 982 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=89430 $Y=11800 $D=1
M1828 999 983 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=89430 $Y=15290 $D=1
M1829 1000 984 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=89430 $Y=18780 $D=1
M1830 1001 985 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=89430 $Y=22270 $D=1
M1831 1002 986 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=89430 $Y=25760 $D=1
M1832 1003 987 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=89430 $Y=29250 $D=1
M1833 1004 988 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=89430 $Y=32740 $D=1
M1834 1005 989 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=89430 $Y=36230 $D=1
M1835 1006 990 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=89430 $Y=39720 $D=1
M1836 1007 991 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=89430 $Y=43210 $D=1
M1837 1008 992 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=89430 $Y=46700 $D=1
M1838 1009 993 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=89430 $Y=50190 $D=1
M1839 1010 994 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=89430 $Y=53680 $D=1
M1840 995 WL15 BL28 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=89870 $Y=1085 $D=1
M1841 996 WL14 BL28 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=89870 $Y=4575 $D=1
M1842 997 WL13 BL28 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=89870 $Y=8065 $D=1
M1843 998 WL12 BL28 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=89870 $Y=11555 $D=1
M1844 999 WL11 BL28 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=89870 $Y=15045 $D=1
M1845 1000 WL10 BL28 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=89870 $Y=18535 $D=1
M1846 1001 WL9 BL28 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=89870 $Y=22025 $D=1
M1847 1002 WL8 BL28 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=89870 $Y=25515 $D=1
M1848 1003 WL7 BL28 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=89870 $Y=29005 $D=1
M1849 1004 WL6 BL28 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=89870 $Y=32495 $D=1
M1850 1005 WL5 BL28 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=89870 $Y=35985 $D=1
M1851 1006 WL4 BL28 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=89870 $Y=39475 $D=1
M1852 1007 WL3 BL28 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=89870 $Y=42965 $D=1
M1853 1008 WL2 BL28 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=89870 $Y=46455 $D=1
M1854 1009 WL1 BL28 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=89870 $Y=49945 $D=1
M1855 1010 WL0 BL28 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=89870 $Y=53435 $D=1
M1856 1011 WL15 !BL29 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=91220 $Y=1085 $D=1
M1857 1012 WL14 !BL29 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=91220 $Y=4575 $D=1
M1858 1013 WL13 !BL29 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=91220 $Y=8065 $D=1
M1859 1014 WL12 !BL29 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=91220 $Y=11555 $D=1
M1860 1015 WL11 !BL29 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=91220 $Y=15045 $D=1
M1861 1016 WL10 !BL29 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=91220 $Y=18535 $D=1
M1862 1017 WL9 !BL29 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=91220 $Y=22025 $D=1
M1863 1018 WL8 !BL29 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=91220 $Y=25515 $D=1
M1864 1019 WL7 !BL29 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=91220 $Y=29005 $D=1
M1865 1020 WL6 !BL29 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=91220 $Y=32495 $D=1
M1866 1021 WL5 !BL29 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=91220 $Y=35985 $D=1
M1867 1022 WL4 !BL29 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=91220 $Y=39475 $D=1
M1868 1023 WL3 !BL29 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=91220 $Y=42965 $D=1
M1869 1024 WL2 !BL29 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=91220 $Y=46455 $D=1
M1870 1025 WL1 !BL29 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=91220 $Y=49945 $D=1
M1871 1026 WL0 !BL29 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=91220 $Y=53435 $D=1
M1872 gnd! 1027 1011 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=91945 $Y=1330 $D=1
M1873 gnd! 1028 1012 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=91945 $Y=4820 $D=1
M1874 gnd! 1029 1013 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=91945 $Y=8310 $D=1
M1875 gnd! 1030 1014 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=91945 $Y=11800 $D=1
M1876 gnd! 1031 1015 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=91945 $Y=15290 $D=1
M1877 gnd! 1032 1016 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=91945 $Y=18780 $D=1
M1878 gnd! 1033 1017 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=91945 $Y=22270 $D=1
M1879 gnd! 1034 1018 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=91945 $Y=25760 $D=1
M1880 gnd! 1035 1019 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=91945 $Y=29250 $D=1
M1881 gnd! 1036 1020 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=91945 $Y=32740 $D=1
M1882 gnd! 1037 1021 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=91945 $Y=36230 $D=1
M1883 gnd! 1038 1022 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=91945 $Y=39720 $D=1
M1884 gnd! 1039 1023 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=91945 $Y=43210 $D=1
M1885 gnd! 1040 1024 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=91945 $Y=46700 $D=1
M1886 gnd! 1041 1025 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=91945 $Y=50190 $D=1
M1887 gnd! 1042 1026 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=91945 $Y=53680 $D=1
M1888 1027 1011 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=92535 $Y=1330 $D=1
M1889 1028 1012 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=92535 $Y=4820 $D=1
M1890 1029 1013 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=92535 $Y=8310 $D=1
M1891 1030 1014 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=92535 $Y=11800 $D=1
M1892 1031 1015 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=92535 $Y=15290 $D=1
M1893 1032 1016 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=92535 $Y=18780 $D=1
M1894 1033 1017 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=92535 $Y=22270 $D=1
M1895 1034 1018 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=92535 $Y=25760 $D=1
M1896 1035 1019 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=92535 $Y=29250 $D=1
M1897 1036 1020 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=92535 $Y=32740 $D=1
M1898 1037 1021 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=92535 $Y=36230 $D=1
M1899 1038 1022 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=92535 $Y=39720 $D=1
M1900 1039 1023 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=92535 $Y=43210 $D=1
M1901 1040 1024 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=92535 $Y=46700 $D=1
M1902 1041 1025 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=92535 $Y=50190 $D=1
M1903 1042 1026 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=92535 $Y=53680 $D=1
M1904 1027 WL15 BL29 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=92975 $Y=1085 $D=1
M1905 1028 WL14 BL29 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=92975 $Y=4575 $D=1
M1906 1029 WL13 BL29 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=92975 $Y=8065 $D=1
M1907 1030 WL12 BL29 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=92975 $Y=11555 $D=1
M1908 1031 WL11 BL29 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=92975 $Y=15045 $D=1
M1909 1032 WL10 BL29 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=92975 $Y=18535 $D=1
M1910 1033 WL9 BL29 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=92975 $Y=22025 $D=1
M1911 1034 WL8 BL29 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=92975 $Y=25515 $D=1
M1912 1035 WL7 BL29 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=92975 $Y=29005 $D=1
M1913 1036 WL6 BL29 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=92975 $Y=32495 $D=1
M1914 1037 WL5 BL29 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=92975 $Y=35985 $D=1
M1915 1038 WL4 BL29 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=92975 $Y=39475 $D=1
M1916 1039 WL3 BL29 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=92975 $Y=42965 $D=1
M1917 1040 WL2 BL29 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=92975 $Y=46455 $D=1
M1918 1041 WL1 BL29 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=92975 $Y=49945 $D=1
M1919 1042 WL0 BL29 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=92975 $Y=53435 $D=1
M1920 1043 WL15 !BL30 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=94325 $Y=1085 $D=1
M1921 1044 WL14 !BL30 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=94325 $Y=4575 $D=1
M1922 1045 WL13 !BL30 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=94325 $Y=8065 $D=1
M1923 1046 WL12 !BL30 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=94325 $Y=11555 $D=1
M1924 1047 WL11 !BL30 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=94325 $Y=15045 $D=1
M1925 1048 WL10 !BL30 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=94325 $Y=18535 $D=1
M1926 1049 WL9 !BL30 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=94325 $Y=22025 $D=1
M1927 1050 WL8 !BL30 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=94325 $Y=25515 $D=1
M1928 1051 WL7 !BL30 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=94325 $Y=29005 $D=1
M1929 1052 WL6 !BL30 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=94325 $Y=32495 $D=1
M1930 1053 WL5 !BL30 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=94325 $Y=35985 $D=1
M1931 1054 WL4 !BL30 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=94325 $Y=39475 $D=1
M1932 1055 WL3 !BL30 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=94325 $Y=42965 $D=1
M1933 1056 WL2 !BL30 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=94325 $Y=46455 $D=1
M1934 1057 WL1 !BL30 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=94325 $Y=49945 $D=1
M1935 1058 WL0 !BL30 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=94325 $Y=53435 $D=1
M1936 gnd! 1059 1043 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=95050 $Y=1330 $D=1
M1937 gnd! 1060 1044 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=95050 $Y=4820 $D=1
M1938 gnd! 1061 1045 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=95050 $Y=8310 $D=1
M1939 gnd! 1062 1046 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=95050 $Y=11800 $D=1
M1940 gnd! 1063 1047 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=95050 $Y=15290 $D=1
M1941 gnd! 1064 1048 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=95050 $Y=18780 $D=1
M1942 gnd! 1065 1049 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=95050 $Y=22270 $D=1
M1943 gnd! 1066 1050 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=95050 $Y=25760 $D=1
M1944 gnd! 1067 1051 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=95050 $Y=29250 $D=1
M1945 gnd! 1068 1052 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=95050 $Y=32740 $D=1
M1946 gnd! 1069 1053 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=95050 $Y=36230 $D=1
M1947 gnd! 1070 1054 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=95050 $Y=39720 $D=1
M1948 gnd! 1071 1055 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=95050 $Y=43210 $D=1
M1949 gnd! 1072 1056 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=95050 $Y=46700 $D=1
M1950 gnd! 1073 1057 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=95050 $Y=50190 $D=1
M1951 gnd! 1074 1058 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=95050 $Y=53680 $D=1
M1952 1059 1043 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=95640 $Y=1330 $D=1
M1953 1060 1044 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=95640 $Y=4820 $D=1
M1954 1061 1045 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=95640 $Y=8310 $D=1
M1955 1062 1046 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=95640 $Y=11800 $D=1
M1956 1063 1047 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=95640 $Y=15290 $D=1
M1957 1064 1048 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=95640 $Y=18780 $D=1
M1958 1065 1049 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=95640 $Y=22270 $D=1
M1959 1066 1050 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=95640 $Y=25760 $D=1
M1960 1067 1051 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=95640 $Y=29250 $D=1
M1961 1068 1052 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=95640 $Y=32740 $D=1
M1962 1069 1053 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=95640 $Y=36230 $D=1
M1963 1070 1054 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=95640 $Y=39720 $D=1
M1964 1071 1055 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=95640 $Y=43210 $D=1
M1965 1072 1056 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=95640 $Y=46700 $D=1
M1966 1073 1057 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=95640 $Y=50190 $D=1
M1967 1074 1058 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=95640 $Y=53680 $D=1
M1968 1059 WL15 BL30 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=96080 $Y=1085 $D=1
M1969 1060 WL14 BL30 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=96080 $Y=4575 $D=1
M1970 1061 WL13 BL30 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=96080 $Y=8065 $D=1
M1971 1062 WL12 BL30 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=96080 $Y=11555 $D=1
M1972 1063 WL11 BL30 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=96080 $Y=15045 $D=1
M1973 1064 WL10 BL30 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=96080 $Y=18535 $D=1
M1974 1065 WL9 BL30 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=96080 $Y=22025 $D=1
M1975 1066 WL8 BL30 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=96080 $Y=25515 $D=1
M1976 1067 WL7 BL30 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=96080 $Y=29005 $D=1
M1977 1068 WL6 BL30 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=96080 $Y=32495 $D=1
M1978 1069 WL5 BL30 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=96080 $Y=35985 $D=1
M1979 1070 WL4 BL30 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=96080 $Y=39475 $D=1
M1980 1071 WL3 BL30 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=96080 $Y=42965 $D=1
M1981 1072 WL2 BL30 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=96080 $Y=46455 $D=1
M1982 1073 WL1 BL30 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=96080 $Y=49945 $D=1
M1983 1074 WL0 BL30 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=96080 $Y=53435 $D=1
M1984 1075 WL15 !BL31 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=97430 $Y=1085 $D=1
M1985 1076 WL14 !BL31 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=97430 $Y=4575 $D=1
M1986 1077 WL13 !BL31 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=97430 $Y=8065 $D=1
M1987 1078 WL12 !BL31 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=97430 $Y=11555 $D=1
M1988 1079 WL11 !BL31 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=97430 $Y=15045 $D=1
M1989 1080 WL10 !BL31 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=97430 $Y=18535 $D=1
M1990 1081 WL9 !BL31 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=97430 $Y=22025 $D=1
M1991 1082 WL8 !BL31 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=97430 $Y=25515 $D=1
M1992 1083 WL7 !BL31 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=97430 $Y=29005 $D=1
M1993 1084 WL6 !BL31 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=97430 $Y=32495 $D=1
M1994 1085 WL5 !BL31 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=97430 $Y=35985 $D=1
M1995 1086 WL4 !BL31 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=97430 $Y=39475 $D=1
M1996 1087 WL3 !BL31 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=97430 $Y=42965 $D=1
M1997 1088 WL2 !BL31 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=97430 $Y=46455 $D=1
M1998 1089 WL1 !BL31 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=97430 $Y=49945 $D=1
M1999 1090 WL0 !BL31 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=97430 $Y=53435 $D=1
M2000 gnd! 1091 1075 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=98155 $Y=1330 $D=1
M2001 gnd! 1092 1076 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=98155 $Y=4820 $D=1
M2002 gnd! 1093 1077 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=98155 $Y=8310 $D=1
M2003 gnd! 1094 1078 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=98155 $Y=11800 $D=1
M2004 gnd! 1095 1079 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=98155 $Y=15290 $D=1
M2005 gnd! 1096 1080 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=98155 $Y=18780 $D=1
M2006 gnd! 1097 1081 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=98155 $Y=22270 $D=1
M2007 gnd! 1098 1082 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=98155 $Y=25760 $D=1
M2008 gnd! 1099 1083 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=98155 $Y=29250 $D=1
M2009 gnd! 1100 1084 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=98155 $Y=32740 $D=1
M2010 gnd! 1101 1085 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=98155 $Y=36230 $D=1
M2011 gnd! 1102 1086 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=98155 $Y=39720 $D=1
M2012 gnd! 1103 1087 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=98155 $Y=43210 $D=1
M2013 gnd! 1104 1088 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=98155 $Y=46700 $D=1
M2014 gnd! 1105 1089 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=98155 $Y=50190 $D=1
M2015 gnd! 1106 1090 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=98155 $Y=53680 $D=1
M2016 1091 1075 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=98745 $Y=1330 $D=1
M2017 1092 1076 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=98745 $Y=4820 $D=1
M2018 1093 1077 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=98745 $Y=8310 $D=1
M2019 1094 1078 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=98745 $Y=11800 $D=1
M2020 1095 1079 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=98745 $Y=15290 $D=1
M2021 1096 1080 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=98745 $Y=18780 $D=1
M2022 1097 1081 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=98745 $Y=22270 $D=1
M2023 1098 1082 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=98745 $Y=25760 $D=1
M2024 1099 1083 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=98745 $Y=29250 $D=1
M2025 1100 1084 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=98745 $Y=32740 $D=1
M2026 1101 1085 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=98745 $Y=36230 $D=1
M2027 1102 1086 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=98745 $Y=39720 $D=1
M2028 1103 1087 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=98745 $Y=43210 $D=1
M2029 1104 1088 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=98745 $Y=46700 $D=1
M2030 1105 1089 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=98745 $Y=50190 $D=1
M2031 1106 1090 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=98745 $Y=53680 $D=1
M2032 1091 WL15 BL31 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=99185 $Y=1085 $D=1
M2033 1092 WL14 BL31 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=99185 $Y=4575 $D=1
M2034 1093 WL13 BL31 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=99185 $Y=8065 $D=1
M2035 1094 WL12 BL31 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=99185 $Y=11555 $D=1
M2036 1095 WL11 BL31 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=99185 $Y=15045 $D=1
M2037 1096 WL10 BL31 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=99185 $Y=18535 $D=1
M2038 1097 WL9 BL31 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=99185 $Y=22025 $D=1
M2039 1098 WL8 BL31 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=99185 $Y=25515 $D=1
M2040 1099 WL7 BL31 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=99185 $Y=29005 $D=1
M2041 1100 WL6 BL31 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=99185 $Y=32495 $D=1
M2042 1101 WL5 BL31 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=99185 $Y=35985 $D=1
M2043 1102 WL4 BL31 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=99185 $Y=39475 $D=1
M2044 1103 WL3 BL31 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=99185 $Y=42965 $D=1
M2045 1104 WL2 BL31 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=99185 $Y=46455 $D=1
M2046 1105 WL1 BL31 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=99185 $Y=49945 $D=1
M2047 1106 WL0 BL31 gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=99185 $Y=53435 $D=1
M2048 BL0 clk vdd! vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=1495 $Y=56355 $D=0
M2049 vdd! 99 82 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=1900 $Y=2775 $D=0
M2050 vdd! 100 83 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=1900 $Y=6265 $D=0
M2051 vdd! 101 84 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=1900 $Y=9755 $D=0
M2052 vdd! 102 85 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=1900 $Y=13245 $D=0
M2053 vdd! 103 86 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=1900 $Y=16735 $D=0
M2054 vdd! 104 87 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=1900 $Y=20225 $D=0
M2055 vdd! 105 88 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=1900 $Y=23715 $D=0
M2056 vdd! 106 89 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=1900 $Y=27205 $D=0
M2057 vdd! 107 90 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=1900 $Y=30695 $D=0
M2058 vdd! 108 91 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=1900 $Y=34185 $D=0
M2059 vdd! 109 92 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=1900 $Y=37675 $D=0
M2060 vdd! 110 93 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=1900 $Y=41165 $D=0
M2061 vdd! 111 94 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=1900 $Y=44655 $D=0
M2062 vdd! 112 95 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=1900 $Y=48145 $D=0
M2063 vdd! 113 96 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=1900 $Y=51635 $D=0
M2064 vdd! 114 97 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=1900 $Y=55125 $D=0
M2065 !BL0 clk BL0 vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=2350 $Y=56355 $D=0
M2066 99 82 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=2490 $Y=2775 $D=0
M2067 100 83 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=2490 $Y=6265 $D=0
M2068 101 84 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=2490 $Y=9755 $D=0
M2069 102 85 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=2490 $Y=13245 $D=0
M2070 103 86 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=2490 $Y=16735 $D=0
M2071 104 87 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=2490 $Y=20225 $D=0
M2072 105 88 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=2490 $Y=23715 $D=0
M2073 106 89 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=2490 $Y=27205 $D=0
M2074 107 90 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=2490 $Y=30695 $D=0
M2075 108 91 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=2490 $Y=34185 $D=0
M2076 109 92 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=2490 $Y=37675 $D=0
M2077 110 93 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=2490 $Y=41165 $D=0
M2078 111 94 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=2490 $Y=44655 $D=0
M2079 112 95 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=2490 $Y=48145 $D=0
M2080 113 96 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=2490 $Y=51635 $D=0
M2081 114 97 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=2490 $Y=55125 $D=0
M2082 vdd! clk !BL0 vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=3215 $Y=56355 $D=0
M2083 BL1 clk vdd! vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=4600 $Y=56355 $D=0
M2084 vdd! 131 115 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=5005 $Y=2775 $D=0
M2085 vdd! 132 116 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=5005 $Y=6265 $D=0
M2086 vdd! 133 117 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=5005 $Y=9755 $D=0
M2087 vdd! 134 118 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=5005 $Y=13245 $D=0
M2088 vdd! 135 119 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=5005 $Y=16735 $D=0
M2089 vdd! 136 120 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=5005 $Y=20225 $D=0
M2090 vdd! 137 121 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=5005 $Y=23715 $D=0
M2091 vdd! 138 122 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=5005 $Y=27205 $D=0
M2092 vdd! 139 123 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=5005 $Y=30695 $D=0
M2093 vdd! 140 124 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=5005 $Y=34185 $D=0
M2094 vdd! 141 125 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=5005 $Y=37675 $D=0
M2095 vdd! 142 126 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=5005 $Y=41165 $D=0
M2096 vdd! 143 127 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=5005 $Y=44655 $D=0
M2097 vdd! 144 128 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=5005 $Y=48145 $D=0
M2098 vdd! 145 129 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=5005 $Y=51635 $D=0
M2099 vdd! 146 130 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=5005 $Y=55125 $D=0
M2100 !BL1 clk BL1 vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=5455 $Y=56355 $D=0
M2101 131 115 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=5595 $Y=2775 $D=0
M2102 132 116 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=5595 $Y=6265 $D=0
M2103 133 117 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=5595 $Y=9755 $D=0
M2104 134 118 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=5595 $Y=13245 $D=0
M2105 135 119 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=5595 $Y=16735 $D=0
M2106 136 120 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=5595 $Y=20225 $D=0
M2107 137 121 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=5595 $Y=23715 $D=0
M2108 138 122 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=5595 $Y=27205 $D=0
M2109 139 123 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=5595 $Y=30695 $D=0
M2110 140 124 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=5595 $Y=34185 $D=0
M2111 141 125 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=5595 $Y=37675 $D=0
M2112 142 126 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=5595 $Y=41165 $D=0
M2113 143 127 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=5595 $Y=44655 $D=0
M2114 144 128 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=5595 $Y=48145 $D=0
M2115 145 129 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=5595 $Y=51635 $D=0
M2116 146 130 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=5595 $Y=55125 $D=0
M2117 vdd! clk !BL1 vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=6320 $Y=56355 $D=0
M2118 BL2 clk vdd! vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=7705 $Y=56355 $D=0
M2119 vdd! 163 147 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=8110 $Y=2775 $D=0
M2120 vdd! 164 148 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=8110 $Y=6265 $D=0
M2121 vdd! 165 149 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=8110 $Y=9755 $D=0
M2122 vdd! 166 150 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=8110 $Y=13245 $D=0
M2123 vdd! 167 151 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=8110 $Y=16735 $D=0
M2124 vdd! 168 152 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=8110 $Y=20225 $D=0
M2125 vdd! 169 153 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=8110 $Y=23715 $D=0
M2126 vdd! 170 154 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=8110 $Y=27205 $D=0
M2127 vdd! 171 155 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=8110 $Y=30695 $D=0
M2128 vdd! 172 156 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=8110 $Y=34185 $D=0
M2129 vdd! 173 157 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=8110 $Y=37675 $D=0
M2130 vdd! 174 158 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=8110 $Y=41165 $D=0
M2131 vdd! 175 159 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=8110 $Y=44655 $D=0
M2132 vdd! 176 160 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=8110 $Y=48145 $D=0
M2133 vdd! 177 161 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=8110 $Y=51635 $D=0
M2134 vdd! 178 162 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=8110 $Y=55125 $D=0
M2135 !BL2 clk BL2 vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=8560 $Y=56355 $D=0
M2136 163 147 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=8700 $Y=2775 $D=0
M2137 164 148 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=8700 $Y=6265 $D=0
M2138 165 149 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=8700 $Y=9755 $D=0
M2139 166 150 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=8700 $Y=13245 $D=0
M2140 167 151 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=8700 $Y=16735 $D=0
M2141 168 152 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=8700 $Y=20225 $D=0
M2142 169 153 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=8700 $Y=23715 $D=0
M2143 170 154 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=8700 $Y=27205 $D=0
M2144 171 155 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=8700 $Y=30695 $D=0
M2145 172 156 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=8700 $Y=34185 $D=0
M2146 173 157 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=8700 $Y=37675 $D=0
M2147 174 158 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=8700 $Y=41165 $D=0
M2148 175 159 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=8700 $Y=44655 $D=0
M2149 176 160 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=8700 $Y=48145 $D=0
M2150 177 161 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=8700 $Y=51635 $D=0
M2151 178 162 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=8700 $Y=55125 $D=0
M2152 vdd! clk !BL2 vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=9425 $Y=56355 $D=0
M2153 BL3 clk vdd! vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=10810 $Y=56355 $D=0
M2154 vdd! 195 179 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=11215 $Y=2775 $D=0
M2155 vdd! 196 180 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=11215 $Y=6265 $D=0
M2156 vdd! 197 181 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=11215 $Y=9755 $D=0
M2157 vdd! 198 182 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=11215 $Y=13245 $D=0
M2158 vdd! 199 183 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=11215 $Y=16735 $D=0
M2159 vdd! 200 184 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=11215 $Y=20225 $D=0
M2160 vdd! 201 185 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=11215 $Y=23715 $D=0
M2161 vdd! 202 186 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=11215 $Y=27205 $D=0
M2162 vdd! 203 187 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=11215 $Y=30695 $D=0
M2163 vdd! 204 188 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=11215 $Y=34185 $D=0
M2164 vdd! 205 189 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=11215 $Y=37675 $D=0
M2165 vdd! 206 190 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=11215 $Y=41165 $D=0
M2166 vdd! 207 191 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=11215 $Y=44655 $D=0
M2167 vdd! 208 192 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=11215 $Y=48145 $D=0
M2168 vdd! 209 193 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=11215 $Y=51635 $D=0
M2169 vdd! 210 194 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=11215 $Y=55125 $D=0
M2170 !BL3 clk BL3 vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=11665 $Y=56355 $D=0
M2171 195 179 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=11805 $Y=2775 $D=0
M2172 196 180 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=11805 $Y=6265 $D=0
M2173 197 181 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=11805 $Y=9755 $D=0
M2174 198 182 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=11805 $Y=13245 $D=0
M2175 199 183 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=11805 $Y=16735 $D=0
M2176 200 184 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=11805 $Y=20225 $D=0
M2177 201 185 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=11805 $Y=23715 $D=0
M2178 202 186 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=11805 $Y=27205 $D=0
M2179 203 187 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=11805 $Y=30695 $D=0
M2180 204 188 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=11805 $Y=34185 $D=0
M2181 205 189 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=11805 $Y=37675 $D=0
M2182 206 190 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=11805 $Y=41165 $D=0
M2183 207 191 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=11805 $Y=44655 $D=0
M2184 208 192 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=11805 $Y=48145 $D=0
M2185 209 193 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=11805 $Y=51635 $D=0
M2186 210 194 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=11805 $Y=55125 $D=0
M2187 vdd! clk !BL3 vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=12530 $Y=56355 $D=0
M2188 BL4 clk vdd! vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=13915 $Y=56355 $D=0
M2189 vdd! 227 211 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=14320 $Y=2775 $D=0
M2190 vdd! 228 212 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=14320 $Y=6265 $D=0
M2191 vdd! 229 213 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=14320 $Y=9755 $D=0
M2192 vdd! 230 214 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=14320 $Y=13245 $D=0
M2193 vdd! 231 215 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=14320 $Y=16735 $D=0
M2194 vdd! 232 216 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=14320 $Y=20225 $D=0
M2195 vdd! 233 217 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=14320 $Y=23715 $D=0
M2196 vdd! 234 218 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=14320 $Y=27205 $D=0
M2197 vdd! 235 219 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=14320 $Y=30695 $D=0
M2198 vdd! 236 220 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=14320 $Y=34185 $D=0
M2199 vdd! 237 221 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=14320 $Y=37675 $D=0
M2200 vdd! 238 222 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=14320 $Y=41165 $D=0
M2201 vdd! 239 223 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=14320 $Y=44655 $D=0
M2202 vdd! 240 224 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=14320 $Y=48145 $D=0
M2203 vdd! 241 225 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=14320 $Y=51635 $D=0
M2204 vdd! 242 226 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=14320 $Y=55125 $D=0
M2205 !BL4 clk BL4 vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=14770 $Y=56355 $D=0
M2206 227 211 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=14910 $Y=2775 $D=0
M2207 228 212 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=14910 $Y=6265 $D=0
M2208 229 213 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=14910 $Y=9755 $D=0
M2209 230 214 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=14910 $Y=13245 $D=0
M2210 231 215 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=14910 $Y=16735 $D=0
M2211 232 216 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=14910 $Y=20225 $D=0
M2212 233 217 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=14910 $Y=23715 $D=0
M2213 234 218 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=14910 $Y=27205 $D=0
M2214 235 219 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=14910 $Y=30695 $D=0
M2215 236 220 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=14910 $Y=34185 $D=0
M2216 237 221 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=14910 $Y=37675 $D=0
M2217 238 222 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=14910 $Y=41165 $D=0
M2218 239 223 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=14910 $Y=44655 $D=0
M2219 240 224 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=14910 $Y=48145 $D=0
M2220 241 225 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=14910 $Y=51635 $D=0
M2221 242 226 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=14910 $Y=55125 $D=0
M2222 vdd! clk !BL4 vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=15635 $Y=56355 $D=0
M2223 BL5 clk vdd! vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=17020 $Y=56355 $D=0
M2224 vdd! 259 243 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=17425 $Y=2775 $D=0
M2225 vdd! 260 244 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=17425 $Y=6265 $D=0
M2226 vdd! 261 245 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=17425 $Y=9755 $D=0
M2227 vdd! 262 246 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=17425 $Y=13245 $D=0
M2228 vdd! 263 247 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=17425 $Y=16735 $D=0
M2229 vdd! 264 248 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=17425 $Y=20225 $D=0
M2230 vdd! 265 249 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=17425 $Y=23715 $D=0
M2231 vdd! 266 250 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=17425 $Y=27205 $D=0
M2232 vdd! 267 251 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=17425 $Y=30695 $D=0
M2233 vdd! 268 252 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=17425 $Y=34185 $D=0
M2234 vdd! 269 253 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=17425 $Y=37675 $D=0
M2235 vdd! 270 254 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=17425 $Y=41165 $D=0
M2236 vdd! 271 255 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=17425 $Y=44655 $D=0
M2237 vdd! 272 256 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=17425 $Y=48145 $D=0
M2238 vdd! 273 257 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=17425 $Y=51635 $D=0
M2239 vdd! 274 258 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=17425 $Y=55125 $D=0
M2240 !BL5 clk BL5 vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=17875 $Y=56355 $D=0
M2241 259 243 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=18015 $Y=2775 $D=0
M2242 260 244 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=18015 $Y=6265 $D=0
M2243 261 245 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=18015 $Y=9755 $D=0
M2244 262 246 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=18015 $Y=13245 $D=0
M2245 263 247 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=18015 $Y=16735 $D=0
M2246 264 248 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=18015 $Y=20225 $D=0
M2247 265 249 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=18015 $Y=23715 $D=0
M2248 266 250 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=18015 $Y=27205 $D=0
M2249 267 251 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=18015 $Y=30695 $D=0
M2250 268 252 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=18015 $Y=34185 $D=0
M2251 269 253 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=18015 $Y=37675 $D=0
M2252 270 254 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=18015 $Y=41165 $D=0
M2253 271 255 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=18015 $Y=44655 $D=0
M2254 272 256 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=18015 $Y=48145 $D=0
M2255 273 257 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=18015 $Y=51635 $D=0
M2256 274 258 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=18015 $Y=55125 $D=0
M2257 vdd! clk !BL5 vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=18740 $Y=56355 $D=0
M2258 BL6 clk vdd! vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=20125 $Y=56355 $D=0
M2259 vdd! 291 275 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=20530 $Y=2775 $D=0
M2260 vdd! 292 276 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=20530 $Y=6265 $D=0
M2261 vdd! 293 277 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=20530 $Y=9755 $D=0
M2262 vdd! 294 278 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=20530 $Y=13245 $D=0
M2263 vdd! 295 279 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=20530 $Y=16735 $D=0
M2264 vdd! 296 280 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=20530 $Y=20225 $D=0
M2265 vdd! 297 281 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=20530 $Y=23715 $D=0
M2266 vdd! 298 282 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=20530 $Y=27205 $D=0
M2267 vdd! 299 283 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=20530 $Y=30695 $D=0
M2268 vdd! 300 284 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=20530 $Y=34185 $D=0
M2269 vdd! 301 285 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=20530 $Y=37675 $D=0
M2270 vdd! 302 286 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=20530 $Y=41165 $D=0
M2271 vdd! 303 287 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=20530 $Y=44655 $D=0
M2272 vdd! 304 288 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=20530 $Y=48145 $D=0
M2273 vdd! 305 289 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=20530 $Y=51635 $D=0
M2274 vdd! 306 290 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=20530 $Y=55125 $D=0
M2275 !BL6 clk BL6 vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=20980 $Y=56355 $D=0
M2276 291 275 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=21120 $Y=2775 $D=0
M2277 292 276 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=21120 $Y=6265 $D=0
M2278 293 277 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=21120 $Y=9755 $D=0
M2279 294 278 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=21120 $Y=13245 $D=0
M2280 295 279 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=21120 $Y=16735 $D=0
M2281 296 280 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=21120 $Y=20225 $D=0
M2282 297 281 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=21120 $Y=23715 $D=0
M2283 298 282 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=21120 $Y=27205 $D=0
M2284 299 283 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=21120 $Y=30695 $D=0
M2285 300 284 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=21120 $Y=34185 $D=0
M2286 301 285 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=21120 $Y=37675 $D=0
M2287 302 286 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=21120 $Y=41165 $D=0
M2288 303 287 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=21120 $Y=44655 $D=0
M2289 304 288 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=21120 $Y=48145 $D=0
M2290 305 289 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=21120 $Y=51635 $D=0
M2291 306 290 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=21120 $Y=55125 $D=0
M2292 vdd! clk !BL6 vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=21845 $Y=56355 $D=0
M2293 BL7 clk vdd! vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=23230 $Y=56355 $D=0
M2294 vdd! 323 307 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=23635 $Y=2775 $D=0
M2295 vdd! 324 308 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=23635 $Y=6265 $D=0
M2296 vdd! 325 309 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=23635 $Y=9755 $D=0
M2297 vdd! 326 310 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=23635 $Y=13245 $D=0
M2298 vdd! 327 311 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=23635 $Y=16735 $D=0
M2299 vdd! 328 312 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=23635 $Y=20225 $D=0
M2300 vdd! 329 313 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=23635 $Y=23715 $D=0
M2301 vdd! 330 314 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=23635 $Y=27205 $D=0
M2302 vdd! 331 315 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=23635 $Y=30695 $D=0
M2303 vdd! 332 316 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=23635 $Y=34185 $D=0
M2304 vdd! 333 317 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=23635 $Y=37675 $D=0
M2305 vdd! 334 318 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=23635 $Y=41165 $D=0
M2306 vdd! 335 319 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=23635 $Y=44655 $D=0
M2307 vdd! 336 320 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=23635 $Y=48145 $D=0
M2308 vdd! 337 321 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=23635 $Y=51635 $D=0
M2309 vdd! 338 322 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=23635 $Y=55125 $D=0
M2310 !BL7 clk BL7 vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=24085 $Y=56355 $D=0
M2311 323 307 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=24225 $Y=2775 $D=0
M2312 324 308 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=24225 $Y=6265 $D=0
M2313 325 309 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=24225 $Y=9755 $D=0
M2314 326 310 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=24225 $Y=13245 $D=0
M2315 327 311 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=24225 $Y=16735 $D=0
M2316 328 312 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=24225 $Y=20225 $D=0
M2317 329 313 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=24225 $Y=23715 $D=0
M2318 330 314 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=24225 $Y=27205 $D=0
M2319 331 315 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=24225 $Y=30695 $D=0
M2320 332 316 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=24225 $Y=34185 $D=0
M2321 333 317 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=24225 $Y=37675 $D=0
M2322 334 318 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=24225 $Y=41165 $D=0
M2323 335 319 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=24225 $Y=44655 $D=0
M2324 336 320 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=24225 $Y=48145 $D=0
M2325 337 321 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=24225 $Y=51635 $D=0
M2326 338 322 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=24225 $Y=55125 $D=0
M2327 vdd! clk !BL7 vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=24950 $Y=56355 $D=0
M2328 BL8 clk vdd! vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=26335 $Y=56355 $D=0
M2329 vdd! 355 339 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=26740 $Y=2775 $D=0
M2330 vdd! 356 340 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=26740 $Y=6265 $D=0
M2331 vdd! 357 341 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=26740 $Y=9755 $D=0
M2332 vdd! 358 342 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=26740 $Y=13245 $D=0
M2333 vdd! 359 343 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=26740 $Y=16735 $D=0
M2334 vdd! 360 344 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=26740 $Y=20225 $D=0
M2335 vdd! 361 345 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=26740 $Y=23715 $D=0
M2336 vdd! 362 346 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=26740 $Y=27205 $D=0
M2337 vdd! 363 347 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=26740 $Y=30695 $D=0
M2338 vdd! 364 348 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=26740 $Y=34185 $D=0
M2339 vdd! 365 349 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=26740 $Y=37675 $D=0
M2340 vdd! 366 350 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=26740 $Y=41165 $D=0
M2341 vdd! 367 351 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=26740 $Y=44655 $D=0
M2342 vdd! 368 352 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=26740 $Y=48145 $D=0
M2343 vdd! 369 353 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=26740 $Y=51635 $D=0
M2344 vdd! 370 354 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=26740 $Y=55125 $D=0
M2345 !BL8 clk BL8 vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=27190 $Y=56355 $D=0
M2346 355 339 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=27330 $Y=2775 $D=0
M2347 356 340 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=27330 $Y=6265 $D=0
M2348 357 341 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=27330 $Y=9755 $D=0
M2349 358 342 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=27330 $Y=13245 $D=0
M2350 359 343 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=27330 $Y=16735 $D=0
M2351 360 344 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=27330 $Y=20225 $D=0
M2352 361 345 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=27330 $Y=23715 $D=0
M2353 362 346 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=27330 $Y=27205 $D=0
M2354 363 347 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=27330 $Y=30695 $D=0
M2355 364 348 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=27330 $Y=34185 $D=0
M2356 365 349 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=27330 $Y=37675 $D=0
M2357 366 350 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=27330 $Y=41165 $D=0
M2358 367 351 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=27330 $Y=44655 $D=0
M2359 368 352 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=27330 $Y=48145 $D=0
M2360 369 353 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=27330 $Y=51635 $D=0
M2361 370 354 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=27330 $Y=55125 $D=0
M2362 vdd! clk !BL8 vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=28055 $Y=56355 $D=0
M2363 BL9 clk vdd! vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=29440 $Y=56355 $D=0
M2364 vdd! 387 371 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=29845 $Y=2775 $D=0
M2365 vdd! 388 372 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=29845 $Y=6265 $D=0
M2366 vdd! 389 373 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=29845 $Y=9755 $D=0
M2367 vdd! 390 374 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=29845 $Y=13245 $D=0
M2368 vdd! 391 375 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=29845 $Y=16735 $D=0
M2369 vdd! 392 376 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=29845 $Y=20225 $D=0
M2370 vdd! 393 377 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=29845 $Y=23715 $D=0
M2371 vdd! 394 378 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=29845 $Y=27205 $D=0
M2372 vdd! 395 379 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=29845 $Y=30695 $D=0
M2373 vdd! 396 380 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=29845 $Y=34185 $D=0
M2374 vdd! 397 381 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=29845 $Y=37675 $D=0
M2375 vdd! 398 382 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=29845 $Y=41165 $D=0
M2376 vdd! 399 383 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=29845 $Y=44655 $D=0
M2377 vdd! 400 384 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=29845 $Y=48145 $D=0
M2378 vdd! 401 385 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=29845 $Y=51635 $D=0
M2379 vdd! 402 386 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=29845 $Y=55125 $D=0
M2380 !BL9 clk BL9 vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=30295 $Y=56355 $D=0
M2381 387 371 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=30435 $Y=2775 $D=0
M2382 388 372 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=30435 $Y=6265 $D=0
M2383 389 373 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=30435 $Y=9755 $D=0
M2384 390 374 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=30435 $Y=13245 $D=0
M2385 391 375 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=30435 $Y=16735 $D=0
M2386 392 376 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=30435 $Y=20225 $D=0
M2387 393 377 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=30435 $Y=23715 $D=0
M2388 394 378 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=30435 $Y=27205 $D=0
M2389 395 379 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=30435 $Y=30695 $D=0
M2390 396 380 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=30435 $Y=34185 $D=0
M2391 397 381 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=30435 $Y=37675 $D=0
M2392 398 382 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=30435 $Y=41165 $D=0
M2393 399 383 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=30435 $Y=44655 $D=0
M2394 400 384 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=30435 $Y=48145 $D=0
M2395 401 385 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=30435 $Y=51635 $D=0
M2396 402 386 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=30435 $Y=55125 $D=0
M2397 vdd! clk !BL9 vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=31160 $Y=56355 $D=0
M2398 BL10 clk vdd! vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=32545 $Y=56355 $D=0
M2399 vdd! 419 403 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=32950 $Y=2775 $D=0
M2400 vdd! 420 404 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=32950 $Y=6265 $D=0
M2401 vdd! 421 405 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=32950 $Y=9755 $D=0
M2402 vdd! 422 406 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=32950 $Y=13245 $D=0
M2403 vdd! 423 407 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=32950 $Y=16735 $D=0
M2404 vdd! 424 408 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=32950 $Y=20225 $D=0
M2405 vdd! 425 409 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=32950 $Y=23715 $D=0
M2406 vdd! 426 410 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=32950 $Y=27205 $D=0
M2407 vdd! 427 411 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=32950 $Y=30695 $D=0
M2408 vdd! 428 412 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=32950 $Y=34185 $D=0
M2409 vdd! 429 413 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=32950 $Y=37675 $D=0
M2410 vdd! 430 414 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=32950 $Y=41165 $D=0
M2411 vdd! 431 415 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=32950 $Y=44655 $D=0
M2412 vdd! 432 416 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=32950 $Y=48145 $D=0
M2413 vdd! 433 417 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=32950 $Y=51635 $D=0
M2414 vdd! 434 418 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=32950 $Y=55125 $D=0
M2415 !BL10 clk BL10 vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=33400 $Y=56355 $D=0
M2416 419 403 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=33540 $Y=2775 $D=0
M2417 420 404 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=33540 $Y=6265 $D=0
M2418 421 405 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=33540 $Y=9755 $D=0
M2419 422 406 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=33540 $Y=13245 $D=0
M2420 423 407 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=33540 $Y=16735 $D=0
M2421 424 408 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=33540 $Y=20225 $D=0
M2422 425 409 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=33540 $Y=23715 $D=0
M2423 426 410 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=33540 $Y=27205 $D=0
M2424 427 411 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=33540 $Y=30695 $D=0
M2425 428 412 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=33540 $Y=34185 $D=0
M2426 429 413 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=33540 $Y=37675 $D=0
M2427 430 414 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=33540 $Y=41165 $D=0
M2428 431 415 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=33540 $Y=44655 $D=0
M2429 432 416 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=33540 $Y=48145 $D=0
M2430 433 417 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=33540 $Y=51635 $D=0
M2431 434 418 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=33540 $Y=55125 $D=0
M2432 vdd! clk !BL10 vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=34265 $Y=56355 $D=0
M2433 BL11 clk vdd! vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=35650 $Y=56355 $D=0
M2434 vdd! 451 435 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=36055 $Y=2775 $D=0
M2435 vdd! 452 436 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=36055 $Y=6265 $D=0
M2436 vdd! 453 437 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=36055 $Y=9755 $D=0
M2437 vdd! 454 438 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=36055 $Y=13245 $D=0
M2438 vdd! 455 439 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=36055 $Y=16735 $D=0
M2439 vdd! 456 440 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=36055 $Y=20225 $D=0
M2440 vdd! 457 441 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=36055 $Y=23715 $D=0
M2441 vdd! 458 442 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=36055 $Y=27205 $D=0
M2442 vdd! 459 443 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=36055 $Y=30695 $D=0
M2443 vdd! 460 444 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=36055 $Y=34185 $D=0
M2444 vdd! 461 445 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=36055 $Y=37675 $D=0
M2445 vdd! 462 446 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=36055 $Y=41165 $D=0
M2446 vdd! 463 447 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=36055 $Y=44655 $D=0
M2447 vdd! 464 448 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=36055 $Y=48145 $D=0
M2448 vdd! 465 449 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=36055 $Y=51635 $D=0
M2449 vdd! 466 450 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=36055 $Y=55125 $D=0
M2450 !BL11 clk BL11 vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=36505 $Y=56355 $D=0
M2451 451 435 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=36645 $Y=2775 $D=0
M2452 452 436 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=36645 $Y=6265 $D=0
M2453 453 437 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=36645 $Y=9755 $D=0
M2454 454 438 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=36645 $Y=13245 $D=0
M2455 455 439 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=36645 $Y=16735 $D=0
M2456 456 440 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=36645 $Y=20225 $D=0
M2457 457 441 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=36645 $Y=23715 $D=0
M2458 458 442 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=36645 $Y=27205 $D=0
M2459 459 443 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=36645 $Y=30695 $D=0
M2460 460 444 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=36645 $Y=34185 $D=0
M2461 461 445 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=36645 $Y=37675 $D=0
M2462 462 446 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=36645 $Y=41165 $D=0
M2463 463 447 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=36645 $Y=44655 $D=0
M2464 464 448 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=36645 $Y=48145 $D=0
M2465 465 449 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=36645 $Y=51635 $D=0
M2466 466 450 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=36645 $Y=55125 $D=0
M2467 vdd! clk !BL11 vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=37370 $Y=56355 $D=0
M2468 BL12 clk vdd! vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=38755 $Y=56355 $D=0
M2469 vdd! 483 467 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=39160 $Y=2775 $D=0
M2470 vdd! 484 468 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=39160 $Y=6265 $D=0
M2471 vdd! 485 469 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=39160 $Y=9755 $D=0
M2472 vdd! 486 470 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=39160 $Y=13245 $D=0
M2473 vdd! 487 471 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=39160 $Y=16735 $D=0
M2474 vdd! 488 472 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=39160 $Y=20225 $D=0
M2475 vdd! 489 473 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=39160 $Y=23715 $D=0
M2476 vdd! 490 474 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=39160 $Y=27205 $D=0
M2477 vdd! 491 475 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=39160 $Y=30695 $D=0
M2478 vdd! 492 476 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=39160 $Y=34185 $D=0
M2479 vdd! 493 477 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=39160 $Y=37675 $D=0
M2480 vdd! 494 478 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=39160 $Y=41165 $D=0
M2481 vdd! 495 479 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=39160 $Y=44655 $D=0
M2482 vdd! 496 480 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=39160 $Y=48145 $D=0
M2483 vdd! 497 481 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=39160 $Y=51635 $D=0
M2484 vdd! 498 482 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=39160 $Y=55125 $D=0
M2485 !BL12 clk BL12 vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=39610 $Y=56355 $D=0
M2486 483 467 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=39750 $Y=2775 $D=0
M2487 484 468 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=39750 $Y=6265 $D=0
M2488 485 469 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=39750 $Y=9755 $D=0
M2489 486 470 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=39750 $Y=13245 $D=0
M2490 487 471 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=39750 $Y=16735 $D=0
M2491 488 472 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=39750 $Y=20225 $D=0
M2492 489 473 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=39750 $Y=23715 $D=0
M2493 490 474 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=39750 $Y=27205 $D=0
M2494 491 475 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=39750 $Y=30695 $D=0
M2495 492 476 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=39750 $Y=34185 $D=0
M2496 493 477 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=39750 $Y=37675 $D=0
M2497 494 478 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=39750 $Y=41165 $D=0
M2498 495 479 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=39750 $Y=44655 $D=0
M2499 496 480 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=39750 $Y=48145 $D=0
M2500 497 481 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=39750 $Y=51635 $D=0
M2501 498 482 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=39750 $Y=55125 $D=0
M2502 vdd! clk !BL12 vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=40475 $Y=56355 $D=0
M2503 BL13 clk vdd! vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=41860 $Y=56355 $D=0
M2504 vdd! 515 499 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=42265 $Y=2775 $D=0
M2505 vdd! 516 500 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=42265 $Y=6265 $D=0
M2506 vdd! 517 501 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=42265 $Y=9755 $D=0
M2507 vdd! 518 502 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=42265 $Y=13245 $D=0
M2508 vdd! 519 503 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=42265 $Y=16735 $D=0
M2509 vdd! 520 504 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=42265 $Y=20225 $D=0
M2510 vdd! 521 505 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=42265 $Y=23715 $D=0
M2511 vdd! 522 506 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=42265 $Y=27205 $D=0
M2512 vdd! 523 507 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=42265 $Y=30695 $D=0
M2513 vdd! 524 508 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=42265 $Y=34185 $D=0
M2514 vdd! 525 509 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=42265 $Y=37675 $D=0
M2515 vdd! 526 510 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=42265 $Y=41165 $D=0
M2516 vdd! 527 511 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=42265 $Y=44655 $D=0
M2517 vdd! 528 512 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=42265 $Y=48145 $D=0
M2518 vdd! 529 513 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=42265 $Y=51635 $D=0
M2519 vdd! 530 514 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=42265 $Y=55125 $D=0
M2520 !BL13 clk BL13 vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=42715 $Y=56355 $D=0
M2521 515 499 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=42855 $Y=2775 $D=0
M2522 516 500 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=42855 $Y=6265 $D=0
M2523 517 501 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=42855 $Y=9755 $D=0
M2524 518 502 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=42855 $Y=13245 $D=0
M2525 519 503 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=42855 $Y=16735 $D=0
M2526 520 504 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=42855 $Y=20225 $D=0
M2527 521 505 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=42855 $Y=23715 $D=0
M2528 522 506 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=42855 $Y=27205 $D=0
M2529 523 507 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=42855 $Y=30695 $D=0
M2530 524 508 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=42855 $Y=34185 $D=0
M2531 525 509 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=42855 $Y=37675 $D=0
M2532 526 510 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=42855 $Y=41165 $D=0
M2533 527 511 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=42855 $Y=44655 $D=0
M2534 528 512 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=42855 $Y=48145 $D=0
M2535 529 513 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=42855 $Y=51635 $D=0
M2536 530 514 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=42855 $Y=55125 $D=0
M2537 vdd! clk !BL13 vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=43580 $Y=56355 $D=0
M2538 BL14 clk vdd! vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=44965 $Y=56355 $D=0
M2539 vdd! 547 531 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=45370 $Y=2775 $D=0
M2540 vdd! 548 532 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=45370 $Y=6265 $D=0
M2541 vdd! 549 533 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=45370 $Y=9755 $D=0
M2542 vdd! 550 534 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=45370 $Y=13245 $D=0
M2543 vdd! 551 535 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=45370 $Y=16735 $D=0
M2544 vdd! 552 536 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=45370 $Y=20225 $D=0
M2545 vdd! 553 537 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=45370 $Y=23715 $D=0
M2546 vdd! 554 538 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=45370 $Y=27205 $D=0
M2547 vdd! 555 539 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=45370 $Y=30695 $D=0
M2548 vdd! 556 540 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=45370 $Y=34185 $D=0
M2549 vdd! 557 541 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=45370 $Y=37675 $D=0
M2550 vdd! 558 542 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=45370 $Y=41165 $D=0
M2551 vdd! 559 543 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=45370 $Y=44655 $D=0
M2552 vdd! 560 544 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=45370 $Y=48145 $D=0
M2553 vdd! 561 545 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=45370 $Y=51635 $D=0
M2554 vdd! 562 546 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=45370 $Y=55125 $D=0
M2555 !BL14 clk BL14 vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=45820 $Y=56355 $D=0
M2556 547 531 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=45960 $Y=2775 $D=0
M2557 548 532 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=45960 $Y=6265 $D=0
M2558 549 533 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=45960 $Y=9755 $D=0
M2559 550 534 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=45960 $Y=13245 $D=0
M2560 551 535 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=45960 $Y=16735 $D=0
M2561 552 536 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=45960 $Y=20225 $D=0
M2562 553 537 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=45960 $Y=23715 $D=0
M2563 554 538 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=45960 $Y=27205 $D=0
M2564 555 539 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=45960 $Y=30695 $D=0
M2565 556 540 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=45960 $Y=34185 $D=0
M2566 557 541 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=45960 $Y=37675 $D=0
M2567 558 542 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=45960 $Y=41165 $D=0
M2568 559 543 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=45960 $Y=44655 $D=0
M2569 560 544 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=45960 $Y=48145 $D=0
M2570 561 545 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=45960 $Y=51635 $D=0
M2571 562 546 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=45960 $Y=55125 $D=0
M2572 vdd! clk !BL14 vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=46685 $Y=56355 $D=0
M2573 BL15 clk vdd! vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=48070 $Y=56355 $D=0
M2574 vdd! 579 563 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=48475 $Y=2775 $D=0
M2575 vdd! 580 564 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=48475 $Y=6265 $D=0
M2576 vdd! 581 565 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=48475 $Y=9755 $D=0
M2577 vdd! 582 566 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=48475 $Y=13245 $D=0
M2578 vdd! 583 567 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=48475 $Y=16735 $D=0
M2579 vdd! 584 568 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=48475 $Y=20225 $D=0
M2580 vdd! 585 569 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=48475 $Y=23715 $D=0
M2581 vdd! 586 570 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=48475 $Y=27205 $D=0
M2582 vdd! 587 571 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=48475 $Y=30695 $D=0
M2583 vdd! 588 572 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=48475 $Y=34185 $D=0
M2584 vdd! 589 573 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=48475 $Y=37675 $D=0
M2585 vdd! 590 574 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=48475 $Y=41165 $D=0
M2586 vdd! 591 575 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=48475 $Y=44655 $D=0
M2587 vdd! 592 576 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=48475 $Y=48145 $D=0
M2588 vdd! 593 577 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=48475 $Y=51635 $D=0
M2589 vdd! 594 578 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=48475 $Y=55125 $D=0
M2590 !BL15 clk BL15 vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=48925 $Y=56355 $D=0
M2591 579 563 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=49065 $Y=2775 $D=0
M2592 580 564 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=49065 $Y=6265 $D=0
M2593 581 565 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=49065 $Y=9755 $D=0
M2594 582 566 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=49065 $Y=13245 $D=0
M2595 583 567 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=49065 $Y=16735 $D=0
M2596 584 568 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=49065 $Y=20225 $D=0
M2597 585 569 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=49065 $Y=23715 $D=0
M2598 586 570 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=49065 $Y=27205 $D=0
M2599 587 571 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=49065 $Y=30695 $D=0
M2600 588 572 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=49065 $Y=34185 $D=0
M2601 589 573 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=49065 $Y=37675 $D=0
M2602 590 574 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=49065 $Y=41165 $D=0
M2603 591 575 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=49065 $Y=44655 $D=0
M2604 592 576 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=49065 $Y=48145 $D=0
M2605 593 577 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=49065 $Y=51635 $D=0
M2606 594 578 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=49065 $Y=55125 $D=0
M2607 vdd! clk !BL15 vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=49790 $Y=56355 $D=0
M2608 BL16 clk vdd! vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=51175 $Y=56355 $D=0
M2609 vdd! 611 595 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=51580 $Y=2775 $D=0
M2610 vdd! 612 596 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=51580 $Y=6265 $D=0
M2611 vdd! 613 597 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=51580 $Y=9755 $D=0
M2612 vdd! 614 598 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=51580 $Y=13245 $D=0
M2613 vdd! 615 599 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=51580 $Y=16735 $D=0
M2614 vdd! 616 600 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=51580 $Y=20225 $D=0
M2615 vdd! 617 601 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=51580 $Y=23715 $D=0
M2616 vdd! 618 602 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=51580 $Y=27205 $D=0
M2617 vdd! 619 603 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=51580 $Y=30695 $D=0
M2618 vdd! 620 604 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=51580 $Y=34185 $D=0
M2619 vdd! 621 605 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=51580 $Y=37675 $D=0
M2620 vdd! 622 606 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=51580 $Y=41165 $D=0
M2621 vdd! 623 607 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=51580 $Y=44655 $D=0
M2622 vdd! 624 608 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=51580 $Y=48145 $D=0
M2623 vdd! 625 609 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=51580 $Y=51635 $D=0
M2624 vdd! 626 610 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=51580 $Y=55125 $D=0
M2625 !BL16 clk BL16 vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=52030 $Y=56355 $D=0
M2626 611 595 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=52170 $Y=2775 $D=0
M2627 612 596 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=52170 $Y=6265 $D=0
M2628 613 597 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=52170 $Y=9755 $D=0
M2629 614 598 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=52170 $Y=13245 $D=0
M2630 615 599 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=52170 $Y=16735 $D=0
M2631 616 600 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=52170 $Y=20225 $D=0
M2632 617 601 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=52170 $Y=23715 $D=0
M2633 618 602 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=52170 $Y=27205 $D=0
M2634 619 603 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=52170 $Y=30695 $D=0
M2635 620 604 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=52170 $Y=34185 $D=0
M2636 621 605 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=52170 $Y=37675 $D=0
M2637 622 606 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=52170 $Y=41165 $D=0
M2638 623 607 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=52170 $Y=44655 $D=0
M2639 624 608 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=52170 $Y=48145 $D=0
M2640 625 609 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=52170 $Y=51635 $D=0
M2641 626 610 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=52170 $Y=55125 $D=0
M2642 vdd! clk !BL16 vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=52895 $Y=56355 $D=0
M2643 BL17 clk vdd! vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=54280 $Y=56355 $D=0
M2644 vdd! 643 627 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=54685 $Y=2775 $D=0
M2645 vdd! 644 628 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=54685 $Y=6265 $D=0
M2646 vdd! 645 629 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=54685 $Y=9755 $D=0
M2647 vdd! 646 630 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=54685 $Y=13245 $D=0
M2648 vdd! 647 631 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=54685 $Y=16735 $D=0
M2649 vdd! 648 632 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=54685 $Y=20225 $D=0
M2650 vdd! 649 633 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=54685 $Y=23715 $D=0
M2651 vdd! 650 634 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=54685 $Y=27205 $D=0
M2652 vdd! 651 635 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=54685 $Y=30695 $D=0
M2653 vdd! 652 636 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=54685 $Y=34185 $D=0
M2654 vdd! 653 637 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=54685 $Y=37675 $D=0
M2655 vdd! 654 638 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=54685 $Y=41165 $D=0
M2656 vdd! 655 639 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=54685 $Y=44655 $D=0
M2657 vdd! 656 640 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=54685 $Y=48145 $D=0
M2658 vdd! 657 641 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=54685 $Y=51635 $D=0
M2659 vdd! 658 642 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=54685 $Y=55125 $D=0
M2660 !BL17 clk BL17 vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=55135 $Y=56355 $D=0
M2661 643 627 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=55275 $Y=2775 $D=0
M2662 644 628 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=55275 $Y=6265 $D=0
M2663 645 629 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=55275 $Y=9755 $D=0
M2664 646 630 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=55275 $Y=13245 $D=0
M2665 647 631 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=55275 $Y=16735 $D=0
M2666 648 632 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=55275 $Y=20225 $D=0
M2667 649 633 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=55275 $Y=23715 $D=0
M2668 650 634 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=55275 $Y=27205 $D=0
M2669 651 635 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=55275 $Y=30695 $D=0
M2670 652 636 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=55275 $Y=34185 $D=0
M2671 653 637 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=55275 $Y=37675 $D=0
M2672 654 638 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=55275 $Y=41165 $D=0
M2673 655 639 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=55275 $Y=44655 $D=0
M2674 656 640 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=55275 $Y=48145 $D=0
M2675 657 641 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=55275 $Y=51635 $D=0
M2676 658 642 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=55275 $Y=55125 $D=0
M2677 vdd! clk !BL17 vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=56000 $Y=56355 $D=0
M2678 BL18 clk vdd! vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=57385 $Y=56355 $D=0
M2679 vdd! 675 659 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=57790 $Y=2775 $D=0
M2680 vdd! 676 660 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=57790 $Y=6265 $D=0
M2681 vdd! 677 661 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=57790 $Y=9755 $D=0
M2682 vdd! 678 662 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=57790 $Y=13245 $D=0
M2683 vdd! 679 663 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=57790 $Y=16735 $D=0
M2684 vdd! 680 664 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=57790 $Y=20225 $D=0
M2685 vdd! 681 665 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=57790 $Y=23715 $D=0
M2686 vdd! 682 666 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=57790 $Y=27205 $D=0
M2687 vdd! 683 667 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=57790 $Y=30695 $D=0
M2688 vdd! 684 668 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=57790 $Y=34185 $D=0
M2689 vdd! 685 669 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=57790 $Y=37675 $D=0
M2690 vdd! 686 670 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=57790 $Y=41165 $D=0
M2691 vdd! 687 671 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=57790 $Y=44655 $D=0
M2692 vdd! 688 672 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=57790 $Y=48145 $D=0
M2693 vdd! 689 673 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=57790 $Y=51635 $D=0
M2694 vdd! 690 674 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=57790 $Y=55125 $D=0
M2695 !BL18 clk BL18 vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=58240 $Y=56355 $D=0
M2696 675 659 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=58380 $Y=2775 $D=0
M2697 676 660 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=58380 $Y=6265 $D=0
M2698 677 661 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=58380 $Y=9755 $D=0
M2699 678 662 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=58380 $Y=13245 $D=0
M2700 679 663 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=58380 $Y=16735 $D=0
M2701 680 664 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=58380 $Y=20225 $D=0
M2702 681 665 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=58380 $Y=23715 $D=0
M2703 682 666 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=58380 $Y=27205 $D=0
M2704 683 667 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=58380 $Y=30695 $D=0
M2705 684 668 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=58380 $Y=34185 $D=0
M2706 685 669 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=58380 $Y=37675 $D=0
M2707 686 670 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=58380 $Y=41165 $D=0
M2708 687 671 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=58380 $Y=44655 $D=0
M2709 688 672 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=58380 $Y=48145 $D=0
M2710 689 673 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=58380 $Y=51635 $D=0
M2711 690 674 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=58380 $Y=55125 $D=0
M2712 vdd! clk !BL18 vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=59105 $Y=56355 $D=0
M2713 BL19 clk vdd! vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=60490 $Y=56355 $D=0
M2714 vdd! 707 691 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=60895 $Y=2775 $D=0
M2715 vdd! 708 692 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=60895 $Y=6265 $D=0
M2716 vdd! 709 693 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=60895 $Y=9755 $D=0
M2717 vdd! 710 694 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=60895 $Y=13245 $D=0
M2718 vdd! 711 695 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=60895 $Y=16735 $D=0
M2719 vdd! 712 696 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=60895 $Y=20225 $D=0
M2720 vdd! 713 697 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=60895 $Y=23715 $D=0
M2721 vdd! 714 698 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=60895 $Y=27205 $D=0
M2722 vdd! 715 699 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=60895 $Y=30695 $D=0
M2723 vdd! 716 700 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=60895 $Y=34185 $D=0
M2724 vdd! 717 701 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=60895 $Y=37675 $D=0
M2725 vdd! 718 702 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=60895 $Y=41165 $D=0
M2726 vdd! 719 703 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=60895 $Y=44655 $D=0
M2727 vdd! 720 704 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=60895 $Y=48145 $D=0
M2728 vdd! 721 705 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=60895 $Y=51635 $D=0
M2729 vdd! 722 706 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=60895 $Y=55125 $D=0
M2730 !BL19 clk BL19 vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=61345 $Y=56355 $D=0
M2731 707 691 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=61485 $Y=2775 $D=0
M2732 708 692 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=61485 $Y=6265 $D=0
M2733 709 693 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=61485 $Y=9755 $D=0
M2734 710 694 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=61485 $Y=13245 $D=0
M2735 711 695 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=61485 $Y=16735 $D=0
M2736 712 696 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=61485 $Y=20225 $D=0
M2737 713 697 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=61485 $Y=23715 $D=0
M2738 714 698 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=61485 $Y=27205 $D=0
M2739 715 699 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=61485 $Y=30695 $D=0
M2740 716 700 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=61485 $Y=34185 $D=0
M2741 717 701 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=61485 $Y=37675 $D=0
M2742 718 702 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=61485 $Y=41165 $D=0
M2743 719 703 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=61485 $Y=44655 $D=0
M2744 720 704 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=61485 $Y=48145 $D=0
M2745 721 705 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=61485 $Y=51635 $D=0
M2746 722 706 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=61485 $Y=55125 $D=0
M2747 vdd! clk !BL19 vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=62210 $Y=56355 $D=0
M2748 BL20 clk vdd! vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=63595 $Y=56355 $D=0
M2749 vdd! 739 723 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=64000 $Y=2775 $D=0
M2750 vdd! 740 724 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=64000 $Y=6265 $D=0
M2751 vdd! 741 725 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=64000 $Y=9755 $D=0
M2752 vdd! 742 726 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=64000 $Y=13245 $D=0
M2753 vdd! 743 727 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=64000 $Y=16735 $D=0
M2754 vdd! 744 728 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=64000 $Y=20225 $D=0
M2755 vdd! 745 729 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=64000 $Y=23715 $D=0
M2756 vdd! 746 730 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=64000 $Y=27205 $D=0
M2757 vdd! 747 731 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=64000 $Y=30695 $D=0
M2758 vdd! 748 732 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=64000 $Y=34185 $D=0
M2759 vdd! 749 733 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=64000 $Y=37675 $D=0
M2760 vdd! 750 734 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=64000 $Y=41165 $D=0
M2761 vdd! 751 735 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=64000 $Y=44655 $D=0
M2762 vdd! 752 736 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=64000 $Y=48145 $D=0
M2763 vdd! 753 737 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=64000 $Y=51635 $D=0
M2764 vdd! 754 738 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=64000 $Y=55125 $D=0
M2765 !BL20 clk BL20 vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=64450 $Y=56355 $D=0
M2766 739 723 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=64590 $Y=2775 $D=0
M2767 740 724 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=64590 $Y=6265 $D=0
M2768 741 725 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=64590 $Y=9755 $D=0
M2769 742 726 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=64590 $Y=13245 $D=0
M2770 743 727 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=64590 $Y=16735 $D=0
M2771 744 728 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=64590 $Y=20225 $D=0
M2772 745 729 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=64590 $Y=23715 $D=0
M2773 746 730 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=64590 $Y=27205 $D=0
M2774 747 731 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=64590 $Y=30695 $D=0
M2775 748 732 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=64590 $Y=34185 $D=0
M2776 749 733 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=64590 $Y=37675 $D=0
M2777 750 734 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=64590 $Y=41165 $D=0
M2778 751 735 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=64590 $Y=44655 $D=0
M2779 752 736 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=64590 $Y=48145 $D=0
M2780 753 737 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=64590 $Y=51635 $D=0
M2781 754 738 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=64590 $Y=55125 $D=0
M2782 vdd! clk !BL20 vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=65315 $Y=56355 $D=0
M2783 BL21 clk vdd! vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=66700 $Y=56355 $D=0
M2784 vdd! 771 755 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=67105 $Y=2775 $D=0
M2785 vdd! 772 756 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=67105 $Y=6265 $D=0
M2786 vdd! 773 757 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=67105 $Y=9755 $D=0
M2787 vdd! 774 758 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=67105 $Y=13245 $D=0
M2788 vdd! 775 759 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=67105 $Y=16735 $D=0
M2789 vdd! 776 760 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=67105 $Y=20225 $D=0
M2790 vdd! 777 761 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=67105 $Y=23715 $D=0
M2791 vdd! 778 762 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=67105 $Y=27205 $D=0
M2792 vdd! 779 763 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=67105 $Y=30695 $D=0
M2793 vdd! 780 764 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=67105 $Y=34185 $D=0
M2794 vdd! 781 765 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=67105 $Y=37675 $D=0
M2795 vdd! 782 766 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=67105 $Y=41165 $D=0
M2796 vdd! 783 767 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=67105 $Y=44655 $D=0
M2797 vdd! 784 768 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=67105 $Y=48145 $D=0
M2798 vdd! 785 769 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=67105 $Y=51635 $D=0
M2799 vdd! 786 770 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=67105 $Y=55125 $D=0
M2800 !BL21 clk BL21 vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=67555 $Y=56355 $D=0
M2801 771 755 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=67695 $Y=2775 $D=0
M2802 772 756 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=67695 $Y=6265 $D=0
M2803 773 757 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=67695 $Y=9755 $D=0
M2804 774 758 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=67695 $Y=13245 $D=0
M2805 775 759 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=67695 $Y=16735 $D=0
M2806 776 760 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=67695 $Y=20225 $D=0
M2807 777 761 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=67695 $Y=23715 $D=0
M2808 778 762 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=67695 $Y=27205 $D=0
M2809 779 763 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=67695 $Y=30695 $D=0
M2810 780 764 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=67695 $Y=34185 $D=0
M2811 781 765 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=67695 $Y=37675 $D=0
M2812 782 766 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=67695 $Y=41165 $D=0
M2813 783 767 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=67695 $Y=44655 $D=0
M2814 784 768 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=67695 $Y=48145 $D=0
M2815 785 769 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=67695 $Y=51635 $D=0
M2816 786 770 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=67695 $Y=55125 $D=0
M2817 vdd! clk !BL21 vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=68420 $Y=56355 $D=0
M2818 BL22 clk vdd! vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=69805 $Y=56355 $D=0
M2819 vdd! 803 787 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=70210 $Y=2775 $D=0
M2820 vdd! 804 788 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=70210 $Y=6265 $D=0
M2821 vdd! 805 789 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=70210 $Y=9755 $D=0
M2822 vdd! 806 790 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=70210 $Y=13245 $D=0
M2823 vdd! 807 791 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=70210 $Y=16735 $D=0
M2824 vdd! 808 792 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=70210 $Y=20225 $D=0
M2825 vdd! 809 793 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=70210 $Y=23715 $D=0
M2826 vdd! 810 794 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=70210 $Y=27205 $D=0
M2827 vdd! 811 795 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=70210 $Y=30695 $D=0
M2828 vdd! 812 796 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=70210 $Y=34185 $D=0
M2829 vdd! 813 797 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=70210 $Y=37675 $D=0
M2830 vdd! 814 798 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=70210 $Y=41165 $D=0
M2831 vdd! 815 799 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=70210 $Y=44655 $D=0
M2832 vdd! 816 800 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=70210 $Y=48145 $D=0
M2833 vdd! 817 801 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=70210 $Y=51635 $D=0
M2834 vdd! 818 802 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=70210 $Y=55125 $D=0
M2835 !BL22 clk BL22 vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=70660 $Y=56355 $D=0
M2836 803 787 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=70800 $Y=2775 $D=0
M2837 804 788 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=70800 $Y=6265 $D=0
M2838 805 789 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=70800 $Y=9755 $D=0
M2839 806 790 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=70800 $Y=13245 $D=0
M2840 807 791 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=70800 $Y=16735 $D=0
M2841 808 792 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=70800 $Y=20225 $D=0
M2842 809 793 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=70800 $Y=23715 $D=0
M2843 810 794 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=70800 $Y=27205 $D=0
M2844 811 795 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=70800 $Y=30695 $D=0
M2845 812 796 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=70800 $Y=34185 $D=0
M2846 813 797 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=70800 $Y=37675 $D=0
M2847 814 798 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=70800 $Y=41165 $D=0
M2848 815 799 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=70800 $Y=44655 $D=0
M2849 816 800 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=70800 $Y=48145 $D=0
M2850 817 801 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=70800 $Y=51635 $D=0
M2851 818 802 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=70800 $Y=55125 $D=0
M2852 vdd! clk !BL22 vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=71525 $Y=56355 $D=0
M2853 BL23 clk vdd! vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=72910 $Y=56355 $D=0
M2854 vdd! 835 819 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=73315 $Y=2775 $D=0
M2855 vdd! 836 820 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=73315 $Y=6265 $D=0
M2856 vdd! 837 821 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=73315 $Y=9755 $D=0
M2857 vdd! 838 822 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=73315 $Y=13245 $D=0
M2858 vdd! 839 823 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=73315 $Y=16735 $D=0
M2859 vdd! 840 824 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=73315 $Y=20225 $D=0
M2860 vdd! 841 825 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=73315 $Y=23715 $D=0
M2861 vdd! 842 826 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=73315 $Y=27205 $D=0
M2862 vdd! 843 827 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=73315 $Y=30695 $D=0
M2863 vdd! 844 828 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=73315 $Y=34185 $D=0
M2864 vdd! 845 829 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=73315 $Y=37675 $D=0
M2865 vdd! 846 830 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=73315 $Y=41165 $D=0
M2866 vdd! 847 831 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=73315 $Y=44655 $D=0
M2867 vdd! 848 832 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=73315 $Y=48145 $D=0
M2868 vdd! 849 833 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=73315 $Y=51635 $D=0
M2869 vdd! 850 834 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=73315 $Y=55125 $D=0
M2870 !BL23 clk BL23 vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=73765 $Y=56355 $D=0
M2871 835 819 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=73905 $Y=2775 $D=0
M2872 836 820 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=73905 $Y=6265 $D=0
M2873 837 821 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=73905 $Y=9755 $D=0
M2874 838 822 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=73905 $Y=13245 $D=0
M2875 839 823 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=73905 $Y=16735 $D=0
M2876 840 824 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=73905 $Y=20225 $D=0
M2877 841 825 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=73905 $Y=23715 $D=0
M2878 842 826 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=73905 $Y=27205 $D=0
M2879 843 827 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=73905 $Y=30695 $D=0
M2880 844 828 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=73905 $Y=34185 $D=0
M2881 845 829 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=73905 $Y=37675 $D=0
M2882 846 830 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=73905 $Y=41165 $D=0
M2883 847 831 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=73905 $Y=44655 $D=0
M2884 848 832 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=73905 $Y=48145 $D=0
M2885 849 833 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=73905 $Y=51635 $D=0
M2886 850 834 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=73905 $Y=55125 $D=0
M2887 vdd! clk !BL23 vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=74630 $Y=56355 $D=0
M2888 BL24 clk vdd! vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=76015 $Y=56355 $D=0
M2889 vdd! 867 851 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=76420 $Y=2775 $D=0
M2890 vdd! 868 852 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=76420 $Y=6265 $D=0
M2891 vdd! 869 853 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=76420 $Y=9755 $D=0
M2892 vdd! 870 854 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=76420 $Y=13245 $D=0
M2893 vdd! 871 855 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=76420 $Y=16735 $D=0
M2894 vdd! 872 856 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=76420 $Y=20225 $D=0
M2895 vdd! 873 857 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=76420 $Y=23715 $D=0
M2896 vdd! 874 858 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=76420 $Y=27205 $D=0
M2897 vdd! 875 859 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=76420 $Y=30695 $D=0
M2898 vdd! 876 860 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=76420 $Y=34185 $D=0
M2899 vdd! 877 861 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=76420 $Y=37675 $D=0
M2900 vdd! 878 862 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=76420 $Y=41165 $D=0
M2901 vdd! 879 863 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=76420 $Y=44655 $D=0
M2902 vdd! 880 864 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=76420 $Y=48145 $D=0
M2903 vdd! 881 865 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=76420 $Y=51635 $D=0
M2904 vdd! 882 866 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=76420 $Y=55125 $D=0
M2905 !BL24 clk BL24 vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=76870 $Y=56355 $D=0
M2906 867 851 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=77010 $Y=2775 $D=0
M2907 868 852 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=77010 $Y=6265 $D=0
M2908 869 853 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=77010 $Y=9755 $D=0
M2909 870 854 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=77010 $Y=13245 $D=0
M2910 871 855 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=77010 $Y=16735 $D=0
M2911 872 856 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=77010 $Y=20225 $D=0
M2912 873 857 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=77010 $Y=23715 $D=0
M2913 874 858 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=77010 $Y=27205 $D=0
M2914 875 859 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=77010 $Y=30695 $D=0
M2915 876 860 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=77010 $Y=34185 $D=0
M2916 877 861 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=77010 $Y=37675 $D=0
M2917 878 862 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=77010 $Y=41165 $D=0
M2918 879 863 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=77010 $Y=44655 $D=0
M2919 880 864 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=77010 $Y=48145 $D=0
M2920 881 865 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=77010 $Y=51635 $D=0
M2921 882 866 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=77010 $Y=55125 $D=0
M2922 vdd! clk !BL24 vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=77735 $Y=56355 $D=0
M2923 BL25 clk vdd! vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=79120 $Y=56355 $D=0
M2924 vdd! 899 883 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=79525 $Y=2775 $D=0
M2925 vdd! 900 884 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=79525 $Y=6265 $D=0
M2926 vdd! 901 885 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=79525 $Y=9755 $D=0
M2927 vdd! 902 886 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=79525 $Y=13245 $D=0
M2928 vdd! 903 887 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=79525 $Y=16735 $D=0
M2929 vdd! 904 888 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=79525 $Y=20225 $D=0
M2930 vdd! 905 889 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=79525 $Y=23715 $D=0
M2931 vdd! 906 890 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=79525 $Y=27205 $D=0
M2932 vdd! 907 891 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=79525 $Y=30695 $D=0
M2933 vdd! 908 892 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=79525 $Y=34185 $D=0
M2934 vdd! 909 893 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=79525 $Y=37675 $D=0
M2935 vdd! 910 894 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=79525 $Y=41165 $D=0
M2936 vdd! 911 895 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=79525 $Y=44655 $D=0
M2937 vdd! 912 896 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=79525 $Y=48145 $D=0
M2938 vdd! 913 897 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=79525 $Y=51635 $D=0
M2939 vdd! 914 898 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=79525 $Y=55125 $D=0
M2940 !BL25 clk BL25 vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=79975 $Y=56355 $D=0
M2941 899 883 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=80115 $Y=2775 $D=0
M2942 900 884 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=80115 $Y=6265 $D=0
M2943 901 885 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=80115 $Y=9755 $D=0
M2944 902 886 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=80115 $Y=13245 $D=0
M2945 903 887 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=80115 $Y=16735 $D=0
M2946 904 888 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=80115 $Y=20225 $D=0
M2947 905 889 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=80115 $Y=23715 $D=0
M2948 906 890 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=80115 $Y=27205 $D=0
M2949 907 891 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=80115 $Y=30695 $D=0
M2950 908 892 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=80115 $Y=34185 $D=0
M2951 909 893 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=80115 $Y=37675 $D=0
M2952 910 894 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=80115 $Y=41165 $D=0
M2953 911 895 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=80115 $Y=44655 $D=0
M2954 912 896 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=80115 $Y=48145 $D=0
M2955 913 897 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=80115 $Y=51635 $D=0
M2956 914 898 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=80115 $Y=55125 $D=0
M2957 vdd! clk !BL25 vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=80840 $Y=56355 $D=0
M2958 BL26 clk vdd! vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=82225 $Y=56355 $D=0
M2959 vdd! 931 915 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=82630 $Y=2775 $D=0
M2960 vdd! 932 916 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=82630 $Y=6265 $D=0
M2961 vdd! 933 917 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=82630 $Y=9755 $D=0
M2962 vdd! 934 918 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=82630 $Y=13245 $D=0
M2963 vdd! 935 919 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=82630 $Y=16735 $D=0
M2964 vdd! 936 920 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=82630 $Y=20225 $D=0
M2965 vdd! 937 921 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=82630 $Y=23715 $D=0
M2966 vdd! 938 922 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=82630 $Y=27205 $D=0
M2967 vdd! 939 923 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=82630 $Y=30695 $D=0
M2968 vdd! 940 924 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=82630 $Y=34185 $D=0
M2969 vdd! 941 925 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=82630 $Y=37675 $D=0
M2970 vdd! 942 926 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=82630 $Y=41165 $D=0
M2971 vdd! 943 927 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=82630 $Y=44655 $D=0
M2972 vdd! 944 928 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=82630 $Y=48145 $D=0
M2973 vdd! 945 929 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=82630 $Y=51635 $D=0
M2974 vdd! 946 930 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=82630 $Y=55125 $D=0
M2975 !BL26 clk BL26 vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=83080 $Y=56355 $D=0
M2976 931 915 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=83220 $Y=2775 $D=0
M2977 932 916 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=83220 $Y=6265 $D=0
M2978 933 917 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=83220 $Y=9755 $D=0
M2979 934 918 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=83220 $Y=13245 $D=0
M2980 935 919 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=83220 $Y=16735 $D=0
M2981 936 920 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=83220 $Y=20225 $D=0
M2982 937 921 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=83220 $Y=23715 $D=0
M2983 938 922 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=83220 $Y=27205 $D=0
M2984 939 923 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=83220 $Y=30695 $D=0
M2985 940 924 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=83220 $Y=34185 $D=0
M2986 941 925 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=83220 $Y=37675 $D=0
M2987 942 926 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=83220 $Y=41165 $D=0
M2988 943 927 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=83220 $Y=44655 $D=0
M2989 944 928 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=83220 $Y=48145 $D=0
M2990 945 929 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=83220 $Y=51635 $D=0
M2991 946 930 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=83220 $Y=55125 $D=0
M2992 vdd! clk !BL26 vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=83945 $Y=56355 $D=0
M2993 BL27 clk vdd! vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=85330 $Y=56355 $D=0
M2994 vdd! 963 947 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=85735 $Y=2775 $D=0
M2995 vdd! 964 948 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=85735 $Y=6265 $D=0
M2996 vdd! 965 949 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=85735 $Y=9755 $D=0
M2997 vdd! 966 950 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=85735 $Y=13245 $D=0
M2998 vdd! 967 951 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=85735 $Y=16735 $D=0
M2999 vdd! 968 952 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=85735 $Y=20225 $D=0
M3000 vdd! 969 953 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=85735 $Y=23715 $D=0
M3001 vdd! 970 954 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=85735 $Y=27205 $D=0
M3002 vdd! 971 955 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=85735 $Y=30695 $D=0
M3003 vdd! 972 956 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=85735 $Y=34185 $D=0
M3004 vdd! 973 957 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=85735 $Y=37675 $D=0
M3005 vdd! 974 958 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=85735 $Y=41165 $D=0
M3006 vdd! 975 959 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=85735 $Y=44655 $D=0
M3007 vdd! 976 960 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=85735 $Y=48145 $D=0
M3008 vdd! 977 961 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=85735 $Y=51635 $D=0
M3009 vdd! 978 962 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=85735 $Y=55125 $D=0
M3010 !BL27 clk BL27 vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=86185 $Y=56355 $D=0
M3011 963 947 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=86325 $Y=2775 $D=0
M3012 964 948 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=86325 $Y=6265 $D=0
M3013 965 949 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=86325 $Y=9755 $D=0
M3014 966 950 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=86325 $Y=13245 $D=0
M3015 967 951 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=86325 $Y=16735 $D=0
M3016 968 952 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=86325 $Y=20225 $D=0
M3017 969 953 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=86325 $Y=23715 $D=0
M3018 970 954 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=86325 $Y=27205 $D=0
M3019 971 955 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=86325 $Y=30695 $D=0
M3020 972 956 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=86325 $Y=34185 $D=0
M3021 973 957 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=86325 $Y=37675 $D=0
M3022 974 958 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=86325 $Y=41165 $D=0
M3023 975 959 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=86325 $Y=44655 $D=0
M3024 976 960 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=86325 $Y=48145 $D=0
M3025 977 961 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=86325 $Y=51635 $D=0
M3026 978 962 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=86325 $Y=55125 $D=0
M3027 vdd! clk !BL27 vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=87050 $Y=56355 $D=0
M3028 BL28 clk vdd! vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=88435 $Y=56355 $D=0
M3029 vdd! 995 979 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=88840 $Y=2775 $D=0
M3030 vdd! 996 980 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=88840 $Y=6265 $D=0
M3031 vdd! 997 981 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=88840 $Y=9755 $D=0
M3032 vdd! 998 982 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=88840 $Y=13245 $D=0
M3033 vdd! 999 983 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=88840 $Y=16735 $D=0
M3034 vdd! 1000 984 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=88840 $Y=20225 $D=0
M3035 vdd! 1001 985 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=88840 $Y=23715 $D=0
M3036 vdd! 1002 986 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=88840 $Y=27205 $D=0
M3037 vdd! 1003 987 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=88840 $Y=30695 $D=0
M3038 vdd! 1004 988 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=88840 $Y=34185 $D=0
M3039 vdd! 1005 989 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=88840 $Y=37675 $D=0
M3040 vdd! 1006 990 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=88840 $Y=41165 $D=0
M3041 vdd! 1007 991 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=88840 $Y=44655 $D=0
M3042 vdd! 1008 992 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=88840 $Y=48145 $D=0
M3043 vdd! 1009 993 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=88840 $Y=51635 $D=0
M3044 vdd! 1010 994 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=88840 $Y=55125 $D=0
M3045 !BL28 clk BL28 vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=89290 $Y=56355 $D=0
M3046 995 979 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=89430 $Y=2775 $D=0
M3047 996 980 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=89430 $Y=6265 $D=0
M3048 997 981 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=89430 $Y=9755 $D=0
M3049 998 982 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=89430 $Y=13245 $D=0
M3050 999 983 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=89430 $Y=16735 $D=0
M3051 1000 984 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=89430 $Y=20225 $D=0
M3052 1001 985 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=89430 $Y=23715 $D=0
M3053 1002 986 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=89430 $Y=27205 $D=0
M3054 1003 987 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=89430 $Y=30695 $D=0
M3055 1004 988 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=89430 $Y=34185 $D=0
M3056 1005 989 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=89430 $Y=37675 $D=0
M3057 1006 990 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=89430 $Y=41165 $D=0
M3058 1007 991 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=89430 $Y=44655 $D=0
M3059 1008 992 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=89430 $Y=48145 $D=0
M3060 1009 993 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=89430 $Y=51635 $D=0
M3061 1010 994 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=89430 $Y=55125 $D=0
M3062 vdd! clk !BL28 vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=90155 $Y=56355 $D=0
M3063 BL29 clk vdd! vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=91540 $Y=56355 $D=0
M3064 vdd! 1027 1011 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=91945 $Y=2775 $D=0
M3065 vdd! 1028 1012 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=91945 $Y=6265 $D=0
M3066 vdd! 1029 1013 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=91945 $Y=9755 $D=0
M3067 vdd! 1030 1014 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=91945 $Y=13245 $D=0
M3068 vdd! 1031 1015 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=91945 $Y=16735 $D=0
M3069 vdd! 1032 1016 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=91945 $Y=20225 $D=0
M3070 vdd! 1033 1017 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=91945 $Y=23715 $D=0
M3071 vdd! 1034 1018 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=91945 $Y=27205 $D=0
M3072 vdd! 1035 1019 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=91945 $Y=30695 $D=0
M3073 vdd! 1036 1020 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=91945 $Y=34185 $D=0
M3074 vdd! 1037 1021 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=91945 $Y=37675 $D=0
M3075 vdd! 1038 1022 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=91945 $Y=41165 $D=0
M3076 vdd! 1039 1023 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=91945 $Y=44655 $D=0
M3077 vdd! 1040 1024 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=91945 $Y=48145 $D=0
M3078 vdd! 1041 1025 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=91945 $Y=51635 $D=0
M3079 vdd! 1042 1026 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=91945 $Y=55125 $D=0
M3080 !BL29 clk BL29 vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=92395 $Y=56355 $D=0
M3081 1027 1011 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=92535 $Y=2775 $D=0
M3082 1028 1012 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=92535 $Y=6265 $D=0
M3083 1029 1013 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=92535 $Y=9755 $D=0
M3084 1030 1014 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=92535 $Y=13245 $D=0
M3085 1031 1015 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=92535 $Y=16735 $D=0
M3086 1032 1016 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=92535 $Y=20225 $D=0
M3087 1033 1017 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=92535 $Y=23715 $D=0
M3088 1034 1018 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=92535 $Y=27205 $D=0
M3089 1035 1019 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=92535 $Y=30695 $D=0
M3090 1036 1020 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=92535 $Y=34185 $D=0
M3091 1037 1021 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=92535 $Y=37675 $D=0
M3092 1038 1022 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=92535 $Y=41165 $D=0
M3093 1039 1023 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=92535 $Y=44655 $D=0
M3094 1040 1024 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=92535 $Y=48145 $D=0
M3095 1041 1025 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=92535 $Y=51635 $D=0
M3096 1042 1026 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=92535 $Y=55125 $D=0
M3097 vdd! clk !BL29 vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=93260 $Y=56355 $D=0
M3098 BL30 clk vdd! vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=94645 $Y=56355 $D=0
M3099 vdd! 1059 1043 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=95050 $Y=2775 $D=0
M3100 vdd! 1060 1044 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=95050 $Y=6265 $D=0
M3101 vdd! 1061 1045 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=95050 $Y=9755 $D=0
M3102 vdd! 1062 1046 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=95050 $Y=13245 $D=0
M3103 vdd! 1063 1047 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=95050 $Y=16735 $D=0
M3104 vdd! 1064 1048 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=95050 $Y=20225 $D=0
M3105 vdd! 1065 1049 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=95050 $Y=23715 $D=0
M3106 vdd! 1066 1050 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=95050 $Y=27205 $D=0
M3107 vdd! 1067 1051 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=95050 $Y=30695 $D=0
M3108 vdd! 1068 1052 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=95050 $Y=34185 $D=0
M3109 vdd! 1069 1053 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=95050 $Y=37675 $D=0
M3110 vdd! 1070 1054 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=95050 $Y=41165 $D=0
M3111 vdd! 1071 1055 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=95050 $Y=44655 $D=0
M3112 vdd! 1072 1056 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=95050 $Y=48145 $D=0
M3113 vdd! 1073 1057 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=95050 $Y=51635 $D=0
M3114 vdd! 1074 1058 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=95050 $Y=55125 $D=0
M3115 !BL30 clk BL30 vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=95500 $Y=56355 $D=0
M3116 1059 1043 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=95640 $Y=2775 $D=0
M3117 1060 1044 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=95640 $Y=6265 $D=0
M3118 1061 1045 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=95640 $Y=9755 $D=0
M3119 1062 1046 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=95640 $Y=13245 $D=0
M3120 1063 1047 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=95640 $Y=16735 $D=0
M3121 1064 1048 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=95640 $Y=20225 $D=0
M3122 1065 1049 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=95640 $Y=23715 $D=0
M3123 1066 1050 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=95640 $Y=27205 $D=0
M3124 1067 1051 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=95640 $Y=30695 $D=0
M3125 1068 1052 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=95640 $Y=34185 $D=0
M3126 1069 1053 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=95640 $Y=37675 $D=0
M3127 1070 1054 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=95640 $Y=41165 $D=0
M3128 1071 1055 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=95640 $Y=44655 $D=0
M3129 1072 1056 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=95640 $Y=48145 $D=0
M3130 1073 1057 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=95640 $Y=51635 $D=0
M3131 1074 1058 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=95640 $Y=55125 $D=0
M3132 vdd! clk !BL30 vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=96365 $Y=56355 $D=0
M3133 BL31 clk vdd! vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=97750 $Y=56355 $D=0
M3134 vdd! 1091 1075 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=98155 $Y=2775 $D=0
M3135 vdd! 1092 1076 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=98155 $Y=6265 $D=0
M3136 vdd! 1093 1077 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=98155 $Y=9755 $D=0
M3137 vdd! 1094 1078 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=98155 $Y=13245 $D=0
M3138 vdd! 1095 1079 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=98155 $Y=16735 $D=0
M3139 vdd! 1096 1080 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=98155 $Y=20225 $D=0
M3140 vdd! 1097 1081 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=98155 $Y=23715 $D=0
M3141 vdd! 1098 1082 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=98155 $Y=27205 $D=0
M3142 vdd! 1099 1083 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=98155 $Y=30695 $D=0
M3143 vdd! 1100 1084 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=98155 $Y=34185 $D=0
M3144 vdd! 1101 1085 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=98155 $Y=37675 $D=0
M3145 vdd! 1102 1086 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=98155 $Y=41165 $D=0
M3146 vdd! 1103 1087 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=98155 $Y=44655 $D=0
M3147 vdd! 1104 1088 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=98155 $Y=48145 $D=0
M3148 vdd! 1105 1089 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=98155 $Y=51635 $D=0
M3149 vdd! 1106 1090 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=98155 $Y=55125 $D=0
M3150 !BL31 clk BL31 vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=98605 $Y=56355 $D=0
M3151 1091 1075 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=98745 $Y=2775 $D=0
M3152 1092 1076 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=98745 $Y=6265 $D=0
M3153 1093 1077 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=98745 $Y=9755 $D=0
M3154 1094 1078 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=98745 $Y=13245 $D=0
M3155 1095 1079 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=98745 $Y=16735 $D=0
M3156 1096 1080 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=98745 $Y=20225 $D=0
M3157 1097 1081 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=98745 $Y=23715 $D=0
M3158 1098 1082 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=98745 $Y=27205 $D=0
M3159 1099 1083 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=98745 $Y=30695 $D=0
M3160 1100 1084 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=98745 $Y=34185 $D=0
M3161 1101 1085 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=98745 $Y=37675 $D=0
M3162 1102 1086 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=98745 $Y=41165 $D=0
M3163 1103 1087 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=98745 $Y=44655 $D=0
M3164 1104 1088 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=98745 $Y=48145 $D=0
M3165 1105 1089 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=98745 $Y=51635 $D=0
M3166 1106 1090 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=98745 $Y=55125 $D=0
M3167 vdd! clk !BL31 vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=99470 $Y=56355 $D=0
.ENDS
***************************************
