* SPICE NETLIST
***************************************

.SUBCKT SRAM_Column gnd! !BL BL WL15 WL14 WL13 WL12 WL11 WL10 WL9 WL8 WL7 WL6 WL5 WL4 WL3 WL2 WL1 WL0 clk
+ vdd!
** N=53 EP=21 IP=0 FDC=99
M0 20 WL15 !BL gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=735 $Y=690 $D=1
M1 21 WL14 !BL gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=735 $Y=4180 $D=1
M2 22 WL13 !BL gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=735 $Y=7670 $D=1
M3 23 WL12 !BL gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=735 $Y=11160 $D=1
M4 24 WL11 !BL gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=735 $Y=14650 $D=1
M5 25 WL10 !BL gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=735 $Y=18140 $D=1
M6 26 WL9 !BL gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=735 $Y=21630 $D=1
M7 27 WL8 !BL gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=735 $Y=25120 $D=1
M8 28 WL7 !BL gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=735 $Y=28610 $D=1
M9 29 WL6 !BL gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=735 $Y=32100 $D=1
M10 30 WL5 !BL gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=735 $Y=35590 $D=1
M11 31 WL4 !BL gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=735 $Y=39080 $D=1
M12 32 WL3 !BL gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=735 $Y=42570 $D=1
M13 33 WL2 !BL gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=735 $Y=46060 $D=1
M14 34 WL1 !BL gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=735 $Y=49550 $D=1
M15 35 WL0 !BL gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.51875e-14 AS=4.1125e-14 PD=1.27e-06 PS=8.2e-07 $X=735 $Y=53040 $D=1
M16 gnd! 37 20 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=1460 $Y=935 $D=1
M17 gnd! 38 21 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=1460 $Y=4425 $D=1
M18 gnd! 39 22 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=1460 $Y=7915 $D=1
M19 gnd! 40 23 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=1460 $Y=11405 $D=1
M20 gnd! 41 24 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=1460 $Y=14895 $D=1
M21 gnd! 42 25 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=1460 $Y=18385 $D=1
M22 gnd! 43 26 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=1460 $Y=21875 $D=1
M23 gnd! 44 27 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=1460 $Y=25365 $D=1
M24 gnd! 45 28 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=1460 $Y=28855 $D=1
M25 gnd! 46 29 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=1460 $Y=32345 $D=1
M26 gnd! 47 30 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=1460 $Y=35835 $D=1
M27 gnd! 48 31 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=1460 $Y=39325 $D=1
M28 gnd! 49 32 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=1460 $Y=42815 $D=1
M29 gnd! 50 33 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=1460 $Y=46305 $D=1
M30 gnd! 51 34 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=1460 $Y=49795 $D=1
M31 gnd! 52 35 gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.65375e-14 AS=8.51875e-14 PD=1.605e-06 PS=1.27e-06 $X=1460 $Y=53285 $D=1
M32 37 20 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=2050 $Y=935 $D=1
M33 38 21 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=2050 $Y=4425 $D=1
M34 39 22 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=2050 $Y=7915 $D=1
M35 40 23 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=2050 $Y=11405 $D=1
M36 41 24 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=2050 $Y=14895 $D=1
M37 42 25 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=2050 $Y=18385 $D=1
M38 43 26 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=2050 $Y=21875 $D=1
M39 44 27 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=2050 $Y=25365 $D=1
M40 45 28 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=2050 $Y=28855 $D=1
M41 46 29 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=2050 $Y=32345 $D=1
M42 47 30 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=2050 $Y=35835 $D=1
M43 48 31 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=2050 $Y=39325 $D=1
M44 49 32 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=2050 $Y=42815 $D=1
M45 50 33 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=2050 $Y=46305 $D=1
M46 51 34 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=2050 $Y=49795 $D=1
M47 52 35 gnd! gnd! NMOS_VTL L=5e-08 W=2e-07 AD=8.16875e-14 AS=8.65375e-14 PD=1.235e-06 PS=1.605e-06 $X=2050 $Y=53285 $D=1
M48 37 WL15 BL gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=2490 $Y=690 $D=1
M49 38 WL14 BL gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=2490 $Y=4180 $D=1
M50 39 WL13 BL gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=2490 $Y=7670 $D=1
M51 40 WL12 BL gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=2490 $Y=11160 $D=1
M52 41 WL11 BL gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=2490 $Y=14650 $D=1
M53 42 WL10 BL gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=2490 $Y=18140 $D=1
M54 43 WL9 BL gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=2490 $Y=21630 $D=1
M55 44 WL8 BL gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=2490 $Y=25120 $D=1
M56 45 WL7 BL gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=2490 $Y=28610 $D=1
M57 46 WL6 BL gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=2490 $Y=32100 $D=1
M58 47 WL5 BL gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=2490 $Y=35590 $D=1
M59 48 WL4 BL gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=2490 $Y=39080 $D=1
M60 49 WL3 BL gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=2490 $Y=42570 $D=1
M61 50 WL2 BL gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=2490 $Y=46060 $D=1
M62 51 WL1 BL gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=2490 $Y=49550 $D=1
M63 52 WL0 BL gnd! NMOS_VTL L=5e-08 W=1.75e-07 AD=8.16875e-14 AS=4.1125e-14 PD=1.235e-06 PS=8.2e-07 $X=2490 $Y=53040 $D=1
M64 BL clk vdd! vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=1055 $Y=55960 $D=0
M65 vdd! 37 20 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=1460 $Y=2380 $D=0
M66 vdd! 38 21 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=1460 $Y=5870 $D=0
M67 vdd! 39 22 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=1460 $Y=9360 $D=0
M68 vdd! 40 23 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=1460 $Y=12850 $D=0
M69 vdd! 41 24 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=1460 $Y=16340 $D=0
M70 vdd! 42 25 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=1460 $Y=19830 $D=0
M71 vdd! 43 26 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=1460 $Y=23320 $D=0
M72 vdd! 44 27 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=1460 $Y=26810 $D=0
M73 vdd! 45 28 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=1460 $Y=30300 $D=0
M74 vdd! 46 29 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=1460 $Y=33790 $D=0
M75 vdd! 47 30 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=1460 $Y=37280 $D=0
M76 vdd! 48 31 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=1460 $Y=40770 $D=0
M77 vdd! 49 32 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=1460 $Y=44260 $D=0
M78 vdd! 50 33 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=1460 $Y=47750 $D=0
M79 vdd! 51 34 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=1460 $Y=51240 $D=0
M80 vdd! 52 35 vdd! PMOS_VTL L=5e-08 W=1e-07 AD=2.45e-14 AS=1.625e-14 PD=6.9e-07 PS=5.25e-07 $X=1460 $Y=54730 $D=0
M81 !BL clk BL vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=1910 $Y=55960 $D=0
M82 37 20 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=2050 $Y=2380 $D=0
M83 38 21 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=2050 $Y=5870 $D=0
M84 39 22 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=2050 $Y=9360 $D=0
M85 40 23 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=2050 $Y=12850 $D=0
M86 41 24 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=2050 $Y=16340 $D=0
M87 42 25 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=2050 $Y=19830 $D=0
M88 43 26 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=2050 $Y=23320 $D=0
M89 44 27 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=2050 $Y=26810 $D=0
M90 45 28 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=2050 $Y=30300 $D=0
M91 46 29 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=2050 $Y=33790 $D=0
M92 47 30 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=2050 $Y=37280 $D=0
M93 48 31 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=2050 $Y=40770 $D=0
M94 49 32 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=2050 $Y=44260 $D=0
M95 50 33 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=2050 $Y=47750 $D=0
M96 51 34 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=2050 $Y=51240 $D=0
M97 52 35 vdd! vdd! PMOS_VTL L=5e-08 W=1e-07 AD=1.725e-14 AS=2.45e-14 PD=5.45e-07 PS=6.9e-07 $X=2050 $Y=54730 $D=0
M98 vdd! clk !BL vdd! PMOS_VTL L=5e-08 W=4e-07 AD=4.1e-14 AS=4.1e-14 PD=1.005e-06 PS=1.005e-06 $X=2775 $Y=55960 $D=0
.ENDS
***************************************
